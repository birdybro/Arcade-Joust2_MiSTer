library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity joust2_bg_sound_bank_a is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of joust2_bg_sound_bank_a is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"D8",X"DD",X"19",X"0A",X"17",X"26",X"0A",X"96",X"16",X"97",X"17",X"0C",X"15",X"26",X"02",X"0C",
		X"14",X"12",X"86",X"14",X"B7",X"20",X"00",X"B6",X"40",X"00",X"C6",X"15",X"F7",X"20",X"01",X"DC",
		X"20",X"2B",X"1F",X"F7",X"60",X"00",X"54",X"4A",X"26",X"13",X"96",X"1F",X"B7",X"78",X"00",X"E6",
		X"A0",X"86",X"08",X"B7",X"78",X"00",X"10",X"9C",X"1D",X"25",X"02",X"86",X"FF",X"DD",X"20",X"F7",
		X"68",X"00",X"DC",X"19",X"3B",X"1A",X"50",X"86",X"34",X"B7",X"40",X"03",X"C6",X"02",X"1F",X"9B",
		X"10",X"CE",X"07",X"FF",X"8E",X"07",X"FF",X"6F",X"84",X"30",X"1F",X"26",X"FA",X"6F",X"84",X"8E",
		X"40",X"00",X"6F",X"03",X"6F",X"02",X"86",X"34",X"A7",X"03",X"86",X"34",X"A7",X"01",X"BD",X"81",
		X"BC",X"BD",X"82",X"01",X"86",X"80",X"97",X"1F",X"97",X"20",X"86",X"14",X"97",X"16",X"97",X"17",
		X"86",X"3C",X"B7",X"40",X"01",X"86",X"3C",X"B7",X"40",X"03",X"8E",X"03",X"E8",X"10",X"83",X"00",
		X"00",X"30",X"1F",X"26",X"F8",X"F6",X"20",X"01",X"2B",X"FB",X"CC",X"30",X"14",X"F7",X"20",X"00",
		X"F6",X"20",X"01",X"2B",X"FB",X"B7",X"20",X"01",X"F6",X"20",X"01",X"2B",X"FB",X"CC",X"FF",X"10",
		X"F7",X"20",X"00",X"F6",X"20",X"01",X"2B",X"FB",X"B7",X"20",X"01",X"F6",X"20",X"01",X"2B",X"FB",
		X"CC",X"01",X"11",X"F7",X"20",X"00",X"F6",X"20",X"01",X"2B",X"FB",X"B7",X"20",X"01",X"F6",X"20",
		X"01",X"2B",X"FB",X"C6",X"14",X"F7",X"20",X"00",X"F6",X"20",X"01",X"2B",X"FB",X"86",X"15",X"B7",
		X"20",X"01",X"86",X"3D",X"B7",X"40",X"01",X"86",X"3D",X"B7",X"40",X"03",X"1C",X"AF",X"8E",X"FF",
		X"FF",X"10",X"83",X"00",X"00",X"10",X"83",X"00",X"00",X"10",X"83",X"00",X"00",X"30",X"1F",X"26",
		X"F0",X"B6",X"40",X"03",X"84",X"FE",X"B7",X"40",X"03",X"1A",X"50",X"C6",X"02",X"8E",X"00",X"00",
		X"86",X"AA",X"A7",X"84",X"A1",X"84",X"26",X"2A",X"A7",X"84",X"A1",X"80",X"26",X"24",X"8C",X"08",
		X"00",X"26",X"EF",X"C6",X"03",X"8E",X"80",X"00",X"4F",X"A0",X"80",X"8C",X"C0",X"00",X"26",X"F9",
		X"81",X"59",X"26",X"0E",X"4F",X"A0",X"80",X"8C",X"00",X"00",X"26",X"F9",X"81",X"55",X"26",X"02",
		X"C6",X"01",X"7F",X"40",X"01",X"86",X"FF",X"B7",X"40",X"00",X"86",X"3C",X"B7",X"40",X"01",X"1F",
		X"98",X"7F",X"40",X"00",X"8E",X"02",X"00",X"30",X"1F",X"26",X"FC",X"7C",X"40",X"00",X"70",X"40",
		X"00",X"8E",X"02",X"00",X"30",X"1F",X"26",X"FC",X"70",X"40",X"00",X"28",X"E7",X"8E",X"01",X"00",
		X"30",X"1F",X"26",X"FC",X"4A",X"26",X"DA",X"8E",X"00",X"00",X"86",X"FF",X"B7",X"40",X"00",X"30",
		X"1F",X"30",X"01",X"30",X"1F",X"26",X"F8",X"8E",X"00",X"00",X"5F",X"E7",X"80",X"8C",X"07",X"FF",
		X"26",X"F9",X"BD",X"81",X"BC",X"BD",X"82",X"01",X"86",X"80",X"97",X"1F",X"97",X"20",X"86",X"14",
		X"97",X"16",X"97",X"17",X"B6",X"40",X"00",X"B6",X"40",X"01",X"8A",X"01",X"B7",X"40",X"01",X"B6",
		X"40",X"03",X"8A",X"01",X"B7",X"40",X"03",X"1C",X"AF",X"7E",X"8A",X"12",X"8E",X"03",X"F9",X"9F",
		X"0E",X"9F",X"10",X"BF",X"03",X"FB",X"CC",X"00",X"00",X"FD",X"03",X"F9",X"86",X"2E",X"8E",X"04",
		X"0C",X"9F",X"12",X"34",X"02",X"1F",X"10",X"C3",X"00",X"13",X"ED",X"84",X"30",X"88",X"13",X"35",
		X"02",X"4A",X"26",X"EF",X"CC",X"00",X"00",X"ED",X"84",X"39",X"B7",X"03",X"F0",X"B6",X"20",X"01",
		X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"B6",X"03",X"F0",X"B7",X"20",X"01",
		X"39",X"86",X"08",X"B7",X"03",X"EF",X"CC",X"02",X"17",X"8E",X"02",X"22",X"C3",X"00",X"18",X"ED",
		X"81",X"7A",X"03",X"EF",X"26",X"F6",X"39",X"6F",X"80",X"83",X"00",X"01",X"26",X"F9",X"39",X"B6",
		X"40",X"03",X"84",X"FE",X"B7",X"40",X"03",X"F6",X"40",X"02",X"C1",X"A2",X"23",X"11",X"10",X"CE",
		X"07",X"FF",X"B6",X"40",X"03",X"8A",X"01",X"B7",X"40",X"03",X"1C",X"AF",X"7E",X"8A",X"12",X"B6",
		X"40",X"03",X"84",X"FE",X"B7",X"40",X"03",X"1A",X"50",X"34",X"04",X"8E",X"87",X"24",X"35",X"04",
		X"4F",X"58",X"89",X"00",X"30",X"8B",X"E6",X"80",X"A6",X"84",X"34",X"02",X"4F",X"58",X"89",X"00",
		X"8E",X"87",X"16",X"AE",X"8B",X"35",X"02",X"6E",X"84",X"10",X"CE",X"07",X"FF",X"BD",X"82",X"9A",
		X"86",X"00",X"8E",X"07",X"FF",X"A7",X"84",X"30",X"1F",X"26",X"FA",X"A7",X"84",X"BD",X"81",X"BC",
		X"BD",X"82",X"01",X"86",X"80",X"97",X"20",X"86",X"14",X"97",X"16",X"97",X"17",X"B6",X"40",X"03",
		X"8A",X"01",X"B7",X"40",X"03",X"1C",X"AF",X"7E",X"8A",X"12",X"34",X"02",X"86",X"20",X"C6",X"E0",
		X"34",X"02",X"86",X"0F",X"BD",X"81",X"EA",X"5C",X"35",X"02",X"4A",X"26",X"F3",X"C6",X"08",X"B6",
		X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"C6",X"07",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",
		X"01",X"5A",X"2A",X"F5",X"35",X"02",X"39",X"10",X"CE",X"07",X"FF",X"34",X"02",X"86",X"0A",X"97",
		X"16",X"20",X"0A",X"10",X"CE",X"07",X"FF",X"34",X"02",X"86",X"14",X"97",X"16",X"BD",X"82",X"01",
		X"7F",X"03",X"E9",X"8E",X"02",X"F2",X"CC",X"00",X"10",X"BD",X"82",X"17",X"35",X"02",X"8E",X"88",
		X"6A",X"48",X"AE",X"86",X"86",X"FF",X"B7",X"03",X"E2",X"B6",X"03",X"E2",X"4C",X"B7",X"03",X"E2",
		X"81",X"08",X"2D",X"03",X"7E",X"83",X"99",X"DE",X"0E",X"EC",X"C4",X"27",X"60",X"E6",X"45",X"C4",
		X"07",X"F1",X"03",X"E2",X"26",X"53",X"A6",X"44",X"2A",X"4F",X"81",X"11",X"27",X"4B",X"34",X"10",
		X"30",X"46",X"CC",X"00",X"0D",X"BD",X"82",X"17",X"35",X"10",X"EC",X"81",X"BF",X"03",X"E5",X"1F",
		X"01",X"A6",X"80",X"A7",X"44",X"AF",X"48",X"BE",X"03",X"E5",X"CC",X"00",X"01",X"ED",X"46",X"DC",
		X"14",X"ED",X"4C",X"EE",X"C4",X"EC",X"C4",X"27",X"B0",X"E6",X"45",X"C4",X"07",X"F1",X"03",X"E2",
		X"26",X"F1",X"A6",X"44",X"2A",X"ED",X"81",X"11",X"27",X"E9",X"BF",X"03",X"E5",X"BD",X"98",X"C2",
		X"BE",X"03",X"E5",X"EC",X"C4",X"27",X"92",X"20",X"E0",X"EE",X"C4",X"20",X"9C",X"BF",X"03",X"E5",
		X"BD",X"98",X"50",X"1F",X"13",X"BE",X"03",X"E5",X"EC",X"81",X"BF",X"03",X"E5",X"1F",X"01",X"A6",
		X"80",X"A7",X"44",X"AF",X"48",X"BE",X"03",X"E5",X"B6",X"03",X"E2",X"A7",X"45",X"CC",X"00",X"01",
		X"ED",X"46",X"DC",X"14",X"ED",X"4C",X"7E",X"82",X"F9",X"B6",X"40",X"03",X"8A",X"01",X"B7",X"40",
		X"03",X"1C",X"AF",X"7E",X"8A",X"12",X"B7",X"03",X"E9",X"10",X"CE",X"07",X"FF",X"B6",X"40",X"03",
		X"8A",X"01",X"B7",X"40",X"03",X"1C",X"AF",X"7E",X"8A",X"12",X"8E",X"88",X"82",X"48",X"AE",X"86",
		X"A6",X"80",X"F6",X"03",X"E3",X"34",X"04",X"B7",X"03",X"E3",X"34",X"02",X"86",X"08",X"B7",X"03",
		X"E2",X"7A",X"03",X"E2",X"2A",X"03",X"7E",X"84",X"9B",X"78",X"03",X"E3",X"24",X"F3",X"34",X"10",
		X"8E",X"03",X"02",X"B6",X"03",X"E2",X"48",X"30",X"86",X"B6",X"03",X"E2",X"C6",X"18",X"3D",X"C3",
		X"03",X"0F",X"ED",X"84",X"8E",X"03",X"D2",X"B6",X"03",X"E2",X"48",X"30",X"86",X"CC",X"00",X"00",
		X"ED",X"84",X"35",X"10",X"DE",X"0E",X"EC",X"C4",X"27",X"63",X"E6",X"45",X"C4",X"07",X"F1",X"03",
		X"E2",X"26",X"56",X"A6",X"44",X"2B",X"52",X"81",X"11",X"27",X"4E",X"34",X"10",X"30",X"46",X"CC",
		X"00",X"0D",X"BD",X"82",X"17",X"35",X"10",X"EC",X"81",X"BF",X"03",X"E5",X"1F",X"01",X"A6",X"80",
		X"84",X"7F",X"A7",X"44",X"AF",X"48",X"BE",X"03",X"E5",X"CC",X"00",X"01",X"ED",X"46",X"DC",X"14",
		X"ED",X"4C",X"EE",X"C4",X"EC",X"C4",X"27",X"89",X"E6",X"45",X"C4",X"07",X"F1",X"03",X"E2",X"26",
		X"F1",X"A6",X"44",X"2B",X"ED",X"81",X"11",X"27",X"E9",X"BF",X"03",X"E5",X"BD",X"98",X"C2",X"BE",
		X"03",X"E5",X"EC",X"C4",X"26",X"E2",X"7E",X"83",X"D1",X"EE",X"C4",X"20",X"99",X"BF",X"03",X"E5",
		X"BD",X"98",X"50",X"1F",X"13",X"BE",X"03",X"E5",X"EC",X"81",X"BF",X"03",X"E5",X"1F",X"01",X"A6",
		X"80",X"84",X"7F",X"A7",X"44",X"AF",X"48",X"BE",X"03",X"E5",X"B6",X"03",X"E2",X"A7",X"45",X"CC",
		X"00",X"01",X"ED",X"46",X"DC",X"14",X"ED",X"4C",X"7E",X"83",X"D1",X"35",X"02",X"B7",X"03",X"E3",
		X"35",X"02",X"BA",X"03",X"E3",X"B7",X"03",X"E3",X"10",X"CE",X"07",X"FF",X"B6",X"40",X"03",X"8A",
		X"01",X"B7",X"40",X"03",X"1C",X"AF",X"7E",X"8A",X"12",X"01",X"02",X"04",X"08",X"10",X"20",X"40",
		X"80",X"8E",X"99",X"1D",X"48",X"EC",X"86",X"34",X"06",X"BE",X"03",X"E7",X"26",X"06",X"BD",X"98",
		X"50",X"BF",X"03",X"E7",X"35",X"06",X"ED",X"08",X"CC",X"00",X"01",X"ED",X"06",X"86",X"11",X"A7",
		X"04",X"86",X"80",X"A7",X"05",X"DC",X"14",X"ED",X"0C",X"86",X"80",X"97",X"20",X"10",X"CE",X"07",
		X"FF",X"B6",X"40",X"03",X"8A",X"01",X"B7",X"40",X"03",X"1C",X"AF",X"7E",X"8A",X"12",X"B7",X"03",
		X"EA",X"B0",X"03",X"EB",X"27",X"27",X"B7",X"03",X"EC",X"B6",X"03",X"EA",X"B7",X"03",X"EB",X"C6",
		X"07",X"34",X"04",X"E6",X"E4",X"8E",X"84",X"B9",X"A6",X"85",X"B5",X"03",X"E3",X"27",X"05",X"BD",
		X"85",X"F2",X"20",X"03",X"BD",X"85",X"3E",X"6A",X"E4",X"2A",X"E8",X"35",X"04",X"10",X"CE",X"07",
		X"FF",X"B6",X"40",X"03",X"8A",X"01",X"B7",X"40",X"03",X"1C",X"AF",X"7E",X"8A",X"12",X"8E",X"01",
		X"00",X"30",X"88",X"20",X"A6",X"85",X"84",X"07",X"B7",X"03",X"EE",X"8E",X"01",X"00",X"CB",X"60",
		X"CB",X"18",X"A6",X"85",X"BB",X"03",X"EC",X"B7",X"03",X"ED",X"B6",X"20",X"01",X"2B",X"FB",X"1A",
		X"50",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"B6",X"03",X"ED",X"B7",X"20",X"01",X"1C",
		X"AF",X"A7",X"85",X"B6",X"03",X"EE",X"85",X"04",X"27",X"77",X"C0",X"08",X"A6",X"85",X"BB",X"03",
		X"EC",X"B7",X"03",X"ED",X"B6",X"20",X"01",X"2B",X"FB",X"1A",X"50",X"F7",X"20",X"00",X"B6",X"20",
		X"01",X"2B",X"FB",X"B6",X"03",X"ED",X"B7",X"20",X"01",X"1C",X"AF",X"A7",X"85",X"B6",X"03",X"EE",
		X"84",X"03",X"27",X"4D",X"C0",X"08",X"A6",X"85",X"BB",X"03",X"EC",X"B7",X"03",X"ED",X"B6",X"20",
		X"01",X"2B",X"FB",X"1A",X"50",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"B6",X"03",X"ED",
		X"B7",X"20",X"01",X"1C",X"AF",X"A7",X"85",X"B6",X"03",X"EE",X"81",X"07",X"26",X"23",X"C0",X"08",
		X"A6",X"85",X"BB",X"03",X"EC",X"B7",X"03",X"ED",X"B6",X"20",X"01",X"2B",X"FB",X"1A",X"50",X"F7",
		X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"B6",X"03",X"ED",X"B7",X"20",X"01",X"1C",X"AF",X"A7",
		X"85",X"39",X"8E",X"01",X"00",X"30",X"88",X"20",X"A6",X"85",X"84",X"07",X"B7",X"03",X"EE",X"8E",
		X"01",X"00",X"CB",X"60",X"CB",X"18",X"A6",X"85",X"BB",X"03",X"EC",X"A7",X"85",X"B6",X"03",X"EE",
		X"85",X"04",X"27",X"29",X"C0",X"08",X"A6",X"85",X"BB",X"03",X"EC",X"A7",X"85",X"B6",X"03",X"EE",
		X"84",X"03",X"27",X"19",X"C0",X"08",X"A6",X"85",X"BB",X"03",X"EC",X"A7",X"85",X"B6",X"03",X"EE",
		X"81",X"07",X"26",X"09",X"C0",X"08",X"A6",X"85",X"BB",X"03",X"EC",X"A7",X"85",X"39",X"86",X"08",
		X"B7",X"03",X"E2",X"7A",X"03",X"E2",X"2A",X"11",X"10",X"CE",X"07",X"FF",X"B6",X"40",X"03",X"8A",
		X"01",X"B7",X"40",X"03",X"1C",X"AF",X"7E",X"8A",X"12",X"78",X"03",X"E3",X"24",X"E5",X"F6",X"03",
		X"E2",X"86",X"04",X"34",X"02",X"CB",X"E0",X"86",X"0F",X"BD",X"81",X"EA",X"CB",X"08",X"6A",X"E4",
		X"26",X"F7",X"35",X"02",X"C6",X"08",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",
		X"B6",X"20",X"01",X"2B",X"FB",X"B6",X"03",X"E2",X"B7",X"20",X"01",X"1C",X"AF",X"C6",X"20",X"FB",
		X"03",X"E2",X"4F",X"1F",X"01",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",
		X"20",X"01",X"2B",X"FB",X"A6",X"89",X"01",X"00",X"B7",X"20",X"01",X"1C",X"AF",X"CB",X"18",X"4F",
		X"1F",X"01",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",
		X"FB",X"A6",X"89",X"01",X"00",X"B7",X"20",X"01",X"1C",X"AF",X"86",X"18",X"B7",X"03",X"E4",X"CB",
		X"08",X"4F",X"1F",X"01",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",
		X"01",X"2B",X"FB",X"A6",X"89",X"01",X"00",X"B7",X"20",X"01",X"1C",X"AF",X"CB",X"08",X"7A",X"03",
		X"E4",X"26",X"DE",X"DE",X"0E",X"EC",X"C4",X"26",X"03",X"7E",X"86",X"43",X"E6",X"45",X"C4",X"07",
		X"F1",X"03",X"E2",X"26",X"0D",X"A6",X"44",X"2B",X"09",X"81",X"11",X"27",X"05",X"BD",X"98",X"C2",
		X"20",X"E3",X"EE",X"C4",X"20",X"DF",X"82",X"69",X"82",X"D3",X"83",X"A6",X"84",X"FE",X"83",X"BA",
		X"86",X"3E",X"84",X"C1",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"02",X"01",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"04",X"01",X"05",X"01",X"06",X"01",X"07",X"01",X"08",X"01",X"09",
		X"01",X"0A",X"01",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"00",X"06",X"01",X"06",X"02",X"06",X"03",X"06",X"04",X"06",X"05",
		X"06",X"06",X"06",X"07",X"06",X"08",X"06",X"09",X"06",X"0A",X"06",X"0B",X"06",X"0A",X"06",X"0D",
		X"06",X"0E",X"06",X"0F",X"02",X"01",X"02",X"02",X"02",X"03",X"02",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"03",X"01",X"03",X"02",X"03",X"04",X"03",X"06",X"03",X"08",
		X"03",X"0A",X"03",X"0C",X"03",X"0E",X"03",X"10",X"03",X"12",X"03",X"16",X"03",X"1E",X"03",X"25",
		X"03",X"30",X"03",X"3B",X"03",X"45",X"03",X"50",X"03",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"04",X"00",X"04",X"01",X"04",X"02",X"04",X"03",X"04",X"04",X"04",X"05",
		X"04",X"06",X"04",X"07",X"06",X"11",X"06",X"12",X"04",X"0A",X"04",X"0B",X"04",X"0C",X"04",X"0D",
		X"04",X"0E",X"04",X"0F",X"04",X"10",X"04",X"11",X"04",X"12",X"04",X"13",X"04",X"14",X"04",X"15",
		X"04",X"16",X"04",X"17",X"04",X"18",X"06",X"13",X"04",X"1A",X"04",X"1B",X"04",X"1C",X"04",X"1D",
		X"04",X"1E",X"04",X"1F",X"04",X"20",X"06",X"10",X"04",X"22",X"AD",X"44",X"BF",X"1E",X"C9",X"8F",
		X"CF",X"97",X"DC",X"21",X"DC",X"4B",X"DC",X"63",X"DC",X"7B",X"DC",X"96",X"DC",X"B4",X"DC",X"CC",
		X"DC",X"E4",X"DC",X"FC",X"DD",X"6F",X"DD",X"F4",X"DE",X"1C",X"DE",X"75",X"DE",X"E2",X"DE",X"FC",
		X"DF",X"16",X"DF",X"27",X"DF",X"68",X"DF",X"E1",X"E0",X"DB",X"E0",X"EE",X"E1",X"01",X"E1",X"1D",
		X"E1",X"7B",X"E1",X"BA",X"E1",X"CD",X"E1",X"E8",X"E2",X"1E",X"E2",X"3A",X"E2",X"4C",X"E2",X"98",
		X"E2",X"C7",X"E3",X"1F",X"E3",X"6B",X"E3",X"C9",X"E4",X"07",X"E4",X"DC",X"E5",X"4C",X"E5",X"CB",
		X"E5",X"F5",X"E6",X"11",X"E6",X"5F",X"E6",X"82",X"89",X"4C",X"89",X"4F",X"89",X"52",X"89",X"55",
		X"89",X"58",X"89",X"5B",X"89",X"5E",X"89",X"61",X"89",X"64",X"89",X"67",X"89",X"6A",X"89",X"6D",
		X"89",X"70",X"89",X"73",X"89",X"76",X"89",X"79",X"89",X"7C",X"89",X"7F",X"89",X"82",X"89",X"85",
		X"89",X"88",X"89",X"8B",X"89",X"8E",X"89",X"91",X"89",X"94",X"89",X"97",X"89",X"9A",X"89",X"9D",
		X"89",X"A0",X"89",X"A3",X"89",X"A6",X"89",X"A9",X"89",X"AC",X"89",X"AF",X"89",X"B2",X"89",X"B5",
		X"89",X"B8",X"89",X"BB",X"89",X"BE",X"89",X"C1",X"89",X"C4",X"89",X"C7",X"89",X"CA",X"89",X"CD",
		X"89",X"D0",X"89",X"D3",X"89",X"D6",X"89",X"D9",X"89",X"DC",X"89",X"DF",X"89",X"E2",X"89",X"E5",
		X"89",X"E8",X"89",X"EB",X"89",X"EE",X"89",X"F1",X"89",X"F4",X"89",X"F7",X"89",X"FA",X"89",X"FD",
		X"8A",X"00",X"8A",X"03",X"8A",X"06",X"8A",X"09",X"8A",X"0C",X"8A",X"0F",X"00",X"08",X"07",X"00",
		X"08",X"78",X"00",X"0F",X"1F",X"00",X"0F",X"80",X"00",X"10",X"FF",X"00",X"11",X"03",X"00",X"12",
		X"FF",X"00",X"12",X"03",X"00",X"14",X"0C",X"00",X"14",X"30",X"00",X"14",X"80",X"00",X"18",X"FF",
		X"00",X"19",X"FF",X"00",X"1B",X"03",X"00",X"1B",X"C0",X"01",X"20",X"07",X"01",X"20",X"38",X"01",
		X"20",X"C0",X"01",X"28",X"7F",X"01",X"30",X"FC",X"01",X"38",X"03",X"01",X"38",X"70",X"01",X"40",
		X"0F",X"01",X"48",X"0F",X"01",X"50",X"0F",X"01",X"58",X"0F",X"01",X"40",X"70",X"01",X"48",X"70",
		X"01",X"50",X"70",X"01",X"58",X"70",X"01",X"60",X"7F",X"01",X"68",X"7F",X"01",X"70",X"7F",X"01",
		X"78",X"7F",X"01",X"80",X"1F",X"01",X"88",X"1F",X"01",X"90",X"1F",X"01",X"98",X"1F",X"01",X"80",
		X"C0",X"01",X"88",X"C0",X"01",X"90",X"C0",X"01",X"98",X"C0",X"01",X"A0",X"1F",X"01",X"A8",X"1F",
		X"01",X"B0",X"1F",X"01",X"B8",X"1F",X"01",X"A0",X"80",X"01",X"A8",X"80",X"01",X"B0",X"80",X"01",
		X"B8",X"80",X"01",X"C0",X"1F",X"01",X"C8",X"1F",X"01",X"D0",X"1F",X"01",X"D8",X"1F",X"01",X"C0",
		X"C0",X"01",X"C8",X"C0",X"01",X"D0",X"C0",X"01",X"D8",X"C0",X"01",X"E0",X"0F",X"01",X"E8",X"0F",
		X"01",X"F0",X"0F",X"01",X"F8",X"0F",X"01",X"E0",X"F0",X"01",X"E8",X"F0",X"01",X"F0",X"F0",X"01",
		X"F8",X"F0",X"B6",X"20",X"01",X"85",X"01",X"27",X"1B",X"B6",X"40",X"00",X"1A",X"50",X"B6",X"20",
		X"01",X"2B",X"FB",X"86",X"14",X"B7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"86",X"15",X"B7",
		X"20",X"01",X"1C",X"AF",X"DE",X"0E",X"EC",X"C4",X"27",X"D8",X"F6",X"40",X"03",X"C4",X"FE",X"F7",
		X"40",X"03",X"EC",X"46",X"1A",X"50",X"93",X"14",X"E3",X"4C",X"9E",X"14",X"AF",X"4C",X"1C",X"AF",
		X"ED",X"46",X"2F",X"0C",X"F6",X"40",X"03",X"CA",X"01",X"F7",X"40",X"03",X"EE",X"C4",X"20",X"D6",
		X"A6",X"44",X"48",X"8E",X"8A",X"84",X"F6",X"40",X"03",X"C4",X"FE",X"F7",X"40",X"03",X"AD",X"96",
		X"34",X"01",X"F6",X"40",X"03",X"CA",X"01",X"F7",X"40",X"03",X"35",X"01",X"2B",X"B8",X"26",X"E0",
		X"EE",X"C4",X"20",X"B2",X"8A",X"B7",X"8B",X"7F",X"8A",X"B4",X"97",X"F6",X"8A",X"B4",X"8A",X"B4",
		X"8A",X"B4",X"8A",X"B4",X"8B",X"E9",X"8F",X"57",X"8F",X"AE",X"8D",X"E5",X"90",X"28",X"90",X"53",
		X"90",X"6F",X"90",X"76",X"90",X"B6",X"97",X"AB",X"90",X"F8",X"91",X"DF",X"92",X"A2",X"93",X"E2",
		X"94",X"D7",X"95",X"C2",X"1C",X"F3",X"39",X"8E",X"84",X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",
		X"B5",X"03",X"E3",X"26",X"14",X"BD",X"8A",X"F9",X"EC",X"46",X"E3",X"81",X"ED",X"46",X"EC",X"81",
		X"E7",X"44",X"AF",X"48",X"1A",X"04",X"1C",X"F7",X"39",X"AE",X"48",X"A6",X"44",X"2B",X"16",X"BD",
		X"8A",X"F9",X"EC",X"46",X"E3",X"81",X"ED",X"46",X"EC",X"81",X"C4",X"7F",X"E7",X"44",X"AF",X"48",
		X"1A",X"04",X"1C",X"F7",X"39",X"30",X"02",X"20",X"CF",X"AE",X"48",X"A6",X"45",X"84",X"07",X"80",
		X"07",X"26",X"17",X"C6",X"0F",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",
		X"20",X"01",X"2B",X"FB",X"4F",X"B7",X"20",X"01",X"1C",X"AF",X"C6",X"08",X"1A",X"50",X"B6",X"20",
		X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"45",X"B7",X"20",X"01",
		X"1C",X"AF",X"C6",X"28",X"EB",X"45",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",
		X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"80",X"B7",X"20",X"01",X"1C",X"AF",X"CB",X"08",X"1A",X"50",
		X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"80",X"B7",
		X"20",X"01",X"1C",X"AF",X"C6",X"08",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",
		X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"45",X"8A",X"78",X"B7",X"20",X"01",X"1C",X"AF",X"39",X"8E",
		X"84",X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",X"B5",X"03",X"E3",X"26",X"2B",X"C6",X"08",X"1A",
		X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"45",
		X"B7",X"20",X"01",X"1C",X"AF",X"AE",X"48",X"EC",X"46",X"E3",X"81",X"ED",X"46",X"A6",X"80",X"A7",
		X"44",X"AF",X"48",X"1A",X"04",X"1C",X"F7",X"39",X"AE",X"48",X"A6",X"44",X"2B",X"E7",X"C6",X"08",
		X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",
		X"45",X"B7",X"20",X"01",X"1C",X"AF",X"EC",X"46",X"E3",X"81",X"ED",X"46",X"A6",X"80",X"84",X"7F",
		X"A7",X"44",X"AF",X"48",X"1A",X"04",X"1C",X"F7",X"39",X"E6",X"45",X"C4",X"07",X"8E",X"84",X"B9",
		X"A6",X"85",X"B5",X"03",X"E3",X"26",X"0F",X"AE",X"48",X"EC",X"81",X"34",X"06",X"A6",X"80",X"A7",
		X"44",X"AF",X"48",X"7E",X"8D",X"18",X"A6",X"44",X"2A",X"64",X"AE",X"48",X"EC",X"81",X"34",X"06",
		X"A6",X"80",X"A7",X"44",X"AF",X"48",X"E6",X"45",X"C4",X"07",X"8E",X"01",X"00",X"30",X"88",X"20",
		X"BF",X"00",X"00",X"AE",X"E1",X"A6",X"80",X"AF",X"E3",X"BE",X"00",X"00",X"30",X"85",X"A7",X"84",
		X"30",X"88",X"18",X"BF",X"00",X"00",X"AE",X"E1",X"A6",X"80",X"AF",X"E3",X"BE",X"00",X"00",X"A7",
		X"84",X"C6",X"18",X"30",X"08",X"BF",X"00",X"00",X"AE",X"E1",X"A6",X"80",X"AF",X"E3",X"BE",X"00",
		X"00",X"A7",X"84",X"30",X"08",X"5A",X"26",X"ED",X"B6",X"03",X"EA",X"27",X"0A",X"B7",X"03",X"EC",
		X"E6",X"45",X"C4",X"07",X"BD",X"85",X"F2",X"35",X"06",X"1A",X"04",X"1C",X"F7",X"39",X"AE",X"48",
		X"EC",X"81",X"34",X"06",X"A6",X"80",X"84",X"7F",X"A7",X"44",X"AF",X"48",X"AE",X"E1",X"C6",X"08",
		X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",
		X"45",X"84",X"07",X"B7",X"20",X"01",X"1C",X"AF",X"C6",X"20",X"EB",X"45",X"4F",X"34",X"06",X"1A",
		X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"80",
		X"B7",X"20",X"01",X"1C",X"AF",X"BF",X"00",X"00",X"AE",X"E1",X"A7",X"84",X"BE",X"00",X"00",X"CB",
		X"18",X"4F",X"34",X"06",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",
		X"01",X"2B",X"FB",X"A6",X"80",X"B7",X"20",X"01",X"1C",X"AF",X"BF",X"00",X"00",X"AE",X"E1",X"A7",
		X"84",X"BE",X"00",X"00",X"86",X"18",X"B7",X"03",X"E4",X"CB",X"08",X"4F",X"34",X"06",X"1A",X"50",
		X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"80",X"B7",
		X"20",X"01",X"1C",X"AF",X"BF",X"00",X"00",X"AE",X"E1",X"A7",X"84",X"BE",X"00",X"00",X"CB",X"08",
		X"7A",X"03",X"E4",X"26",X"D6",X"1C",X"F3",X"39",X"AE",X"E1",X"C6",X"08",X"1A",X"50",X"B6",X"20",
		X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"45",X"84",X"07",X"B7",
		X"20",X"01",X"1C",X"AF",X"C6",X"20",X"EB",X"45",X"4F",X"34",X"06",X"A6",X"84",X"BF",X"00",X"00",
		X"AE",X"E1",X"A7",X"89",X"01",X"00",X"BE",X"00",X"00",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",
		X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"80",X"84",X"3F",X"B7",X"20",X"01",X"1C",
		X"AF",X"CB",X"18",X"4F",X"34",X"06",X"A6",X"84",X"BF",X"00",X"00",X"AE",X"E1",X"A7",X"89",X"01",
		X"00",X"BE",X"00",X"00",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",
		X"01",X"2B",X"FB",X"A6",X"80",X"B7",X"20",X"01",X"1C",X"AF",X"86",X"18",X"B7",X"03",X"E4",X"C6",
		X"40",X"EB",X"45",X"4F",X"34",X"06",X"A6",X"84",X"BF",X"00",X"00",X"AE",X"E1",X"A7",X"89",X"01",
		X"00",X"BE",X"00",X"00",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",
		X"01",X"2B",X"FB",X"A6",X"80",X"B7",X"20",X"01",X"1C",X"AF",X"CB",X"08",X"7A",X"03",X"E4",X"26",
		X"D2",X"C6",X"20",X"EB",X"45",X"4F",X"1F",X"01",X"A6",X"89",X"01",X"00",X"1A",X"50",X"BD",X"81",
		X"EA",X"1C",X"AF",X"B6",X"03",X"EA",X"27",X"0A",X"B7",X"03",X"EC",X"E6",X"45",X"C4",X"07",X"BD",
		X"85",X"3E",X"1C",X"F3",X"39",X"8E",X"84",X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",X"B5",X"03",
		X"E3",X"26",X"03",X"7E",X"8E",X"78",X"A6",X"44",X"2A",X"6C",X"AE",X"48",X"EC",X"81",X"B7",X"03",
		X"EC",X"E7",X"44",X"AF",X"48",X"8E",X"00",X"20",X"30",X"89",X"01",X"00",X"E6",X"45",X"C4",X"07",
		X"30",X"85",X"A6",X"84",X"84",X"07",X"B7",X"03",X"EE",X"30",X"88",X"58",X"A6",X"84",X"BB",X"03",
		X"EC",X"2A",X"02",X"86",X"7F",X"A7",X"84",X"B6",X"03",X"EE",X"85",X"04",X"27",X"35",X"30",X"18",
		X"A6",X"84",X"BB",X"03",X"EC",X"2A",X"02",X"86",X"7F",X"A7",X"84",X"B6",X"03",X"EE",X"84",X"07",
		X"27",X"21",X"30",X"18",X"A6",X"84",X"BB",X"03",X"EC",X"2A",X"02",X"86",X"7F",X"A7",X"84",X"B6",
		X"03",X"EE",X"81",X"03",X"26",X"0D",X"30",X"18",X"A6",X"84",X"BB",X"03",X"EC",X"2A",X"02",X"86",
		X"7F",X"A7",X"84",X"1C",X"F3",X"39",X"AE",X"48",X"EC",X"81",X"B7",X"03",X"EC",X"C4",X"7F",X"E7",
		X"44",X"AF",X"48",X"8E",X"00",X"20",X"20",X"12",X"AE",X"48",X"EC",X"81",X"B7",X"03",X"EC",X"E7",
		X"44",X"AF",X"48",X"8E",X"00",X"20",X"30",X"89",X"01",X"00",X"E6",X"45",X"C4",X"07",X"30",X"85",
		X"A6",X"84",X"84",X"07",X"B7",X"03",X"EE",X"30",X"88",X"58",X"A6",X"84",X"BB",X"03",X"EC",X"2A",
		X"02",X"86",X"7F",X"B7",X"03",X"ED",X"A7",X"84",X"1F",X"10",X"1A",X"50",X"B6",X"20",X"01",X"2B",
		X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"B6",X"03",X"ED",X"B7",X"20",X"01",X"1C",
		X"AF",X"B6",X"03",X"EE",X"85",X"04",X"26",X"03",X"7E",X"8F",X"54",X"30",X"18",X"A6",X"84",X"BB",
		X"03",X"EC",X"2A",X"02",X"86",X"7F",X"B7",X"03",X"ED",X"A7",X"84",X"1F",X"10",X"1A",X"50",X"B6",
		X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"B6",X"03",X"ED",X"B7",
		X"20",X"01",X"1C",X"AF",X"B6",X"03",X"EE",X"84",X"07",X"27",X"59",X"30",X"18",X"A6",X"84",X"BB",
		X"03",X"EC",X"2A",X"02",X"86",X"7F",X"B7",X"03",X"ED",X"A7",X"84",X"1F",X"10",X"1A",X"50",X"B6",
		X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"B6",X"03",X"ED",X"B7",
		X"20",X"01",X"1C",X"AF",X"B6",X"03",X"EE",X"81",X"03",X"26",X"29",X"30",X"18",X"A6",X"84",X"BB",
		X"03",X"EC",X"2A",X"02",X"86",X"7F",X"B7",X"03",X"ED",X"A7",X"84",X"1F",X"10",X"1A",X"50",X"B6",
		X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"B6",X"03",X"ED",X"B7",
		X"20",X"01",X"1C",X"AF",X"1C",X"F3",X"39",X"8E",X"84",X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",
		X"B5",X"03",X"E3",X"27",X"1B",X"A6",X"44",X"2B",X"17",X"AE",X"48",X"A6",X"80",X"34",X"02",X"EC",
		X"81",X"34",X"06",X"A6",X"80",X"84",X"7F",X"A7",X"44",X"AF",X"48",X"8E",X"03",X"02",X"20",X"13",
		X"AE",X"48",X"A6",X"80",X"34",X"02",X"EC",X"81",X"34",X"06",X"A6",X"80",X"A7",X"44",X"AF",X"48",
		X"8E",X"02",X"22",X"E6",X"45",X"C4",X"07",X"58",X"30",X"85",X"EC",X"84",X"C3",X"00",X"03",X"ED",
		X"84",X"1F",X"01",X"35",X"06",X"ED",X"01",X"35",X"02",X"A7",X"84",X"1C",X"F3",X"39",X"8E",X"84",
		X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",X"B5",X"03",X"E3",X"27",X"3A",X"A6",X"44",X"2B",X"36",
		X"8E",X"03",X"02",X"E6",X"45",X"C4",X"07",X"58",X"30",X"85",X"A6",X"94",X"27",X"19",X"4A",X"A7",
		X"94",X"26",X"14",X"EC",X"84",X"83",X"00",X"03",X"ED",X"84",X"AE",X"48",X"A6",X"80",X"84",X"7F",
		X"A7",X"44",X"AF",X"48",X"1C",X"F3",X"39",X"AE",X"84",X"AE",X"01",X"A6",X"80",X"84",X"7F",X"A7",
		X"44",X"AF",X"48",X"1C",X"F3",X"39",X"8E",X"02",X"22",X"E6",X"45",X"C4",X"07",X"58",X"30",X"85",
		X"A6",X"94",X"27",X"17",X"4A",X"A7",X"94",X"26",X"12",X"EC",X"84",X"83",X"00",X"03",X"ED",X"84",
		X"AE",X"48",X"A6",X"80",X"A7",X"44",X"AF",X"48",X"1C",X"F3",X"39",X"AE",X"84",X"AE",X"01",X"A6",
		X"80",X"A7",X"44",X"AF",X"48",X"1C",X"F3",X"39",X"AE",X"48",X"EC",X"81",X"AF",X"48",X"7D",X"03",
		X"E9",X"27",X"15",X"8E",X"98",X"24",X"48",X"AE",X"86",X"58",X"AE",X"85",X"B6",X"03",X"E9",X"4A",
		X"E6",X"86",X"7F",X"03",X"E9",X"7E",X"82",X"3F",X"AE",X"48",X"A6",X"80",X"A7",X"44",X"AF",X"48",
		X"1C",X"F3",X"39",X"AE",X"48",X"A6",X"80",X"A7",X"44",X"AF",X"48",X"F6",X"03",X"E9",X"27",X"0C",
		X"7F",X"03",X"E9",X"5A",X"8E",X"98",X"50",X"E6",X"85",X"7E",X"82",X"3F",X"1C",X"F3",X"39",X"AE",
		X"48",X"E6",X"80",X"7E",X"82",X"3F",X"A6",X"44",X"2B",X"1F",X"8E",X"03",X"D2",X"E6",X"45",X"C4",
		X"07",X"58",X"30",X"85",X"34",X"10",X"AE",X"48",X"EC",X"81",X"AF",X"F1",X"1F",X"01",X"A6",X"80",
		X"84",X"7F",X"A7",X"44",X"AF",X"48",X"1C",X"F3",X"39",X"8E",X"02",X"F2",X"E6",X"45",X"C4",X"07",
		X"58",X"30",X"85",X"34",X"10",X"AE",X"48",X"EC",X"81",X"AF",X"F1",X"1F",X"01",X"A6",X"80",X"A7",
		X"44",X"AF",X"48",X"1C",X"F3",X"39",X"A6",X"44",X"2B",X"05",X"8E",X"03",X"D2",X"20",X"03",X"8E",
		X"02",X"F2",X"E6",X"45",X"C4",X"07",X"58",X"30",X"85",X"34",X"10",X"EC",X"84",X"27",X"16",X"1F",
		X"01",X"A6",X"80",X"E6",X"44",X"2B",X"02",X"84",X"7F",X"A7",X"44",X"AF",X"48",X"CC",X"00",X"00",
		X"ED",X"F1",X"1C",X"F3",X"39",X"AE",X"48",X"A6",X"80",X"E6",X"44",X"2B",X"02",X"84",X"7F",X"A7",
		X"44",X"AF",X"48",X"32",X"62",X"1C",X"F3",X"39",X"E6",X"45",X"C4",X"07",X"8E",X"84",X"B9",X"A6",
		X"85",X"43",X"B4",X"03",X"E3",X"B7",X"03",X"E3",X"86",X"04",X"34",X"02",X"CB",X"E0",X"1A",X"50",
		X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"86",X"0F",X"B7",
		X"20",X"01",X"CB",X"08",X"6A",X"E4",X"26",X"E8",X"35",X"02",X"C6",X"08",X"1A",X"50",X"B6",X"20",
		X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"45",X"84",X"07",X"B7",
		X"20",X"01",X"1C",X"AF",X"C6",X"20",X"EB",X"45",X"4F",X"1F",X"01",X"1A",X"50",X"B6",X"20",X"01",
		X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"89",X"01",X"00",X"B7",X"20",
		X"01",X"1C",X"AF",X"CB",X"18",X"4F",X"1F",X"01",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",
		X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"89",X"01",X"00",X"B7",X"20",X"01",X"1C",X"AF",
		X"86",X"18",X"B7",X"03",X"E4",X"CB",X"08",X"4F",X"1F",X"01",X"1A",X"50",X"B6",X"20",X"01",X"2B",
		X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"89",X"01",X"00",X"B7",X"20",X"01",
		X"1C",X"AF",X"CB",X"08",X"7A",X"03",X"E4",X"26",X"DE",X"34",X"40",X"A6",X"45",X"84",X"07",X"B7",
		X"03",X"E2",X"DE",X"0E",X"EC",X"C4",X"27",X"1F",X"11",X"A3",X"E4",X"27",X"16",X"A6",X"45",X"84",
		X"07",X"B1",X"03",X"E2",X"26",X"0D",X"A6",X"44",X"2B",X"09",X"81",X"11",X"27",X"05",X"BD",X"98",
		X"C2",X"20",X"E1",X"EE",X"C4",X"20",X"DD",X"35",X"40",X"BD",X"98",X"C2",X"1A",X"08",X"39",X"8E",
		X"84",X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",X"B5",X"03",X"E3",X"26",X"14",X"BD",X"92",X"21",
		X"EC",X"46",X"E3",X"81",X"ED",X"46",X"EC",X"81",X"E7",X"44",X"AF",X"48",X"1A",X"04",X"1C",X"F7",
		X"39",X"AE",X"48",X"A6",X"44",X"2B",X"16",X"BD",X"92",X"21",X"EC",X"46",X"E3",X"81",X"ED",X"46",
		X"EC",X"81",X"C4",X"7F",X"E7",X"44",X"AF",X"48",X"1A",X"04",X"1C",X"F7",X"39",X"30",X"03",X"20",
		X"CF",X"AE",X"48",X"C6",X"08",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",
		X"20",X"01",X"2B",X"FB",X"A6",X"45",X"B7",X"20",X"01",X"1C",X"AF",X"C6",X"0F",X"1A",X"50",X"B6",
		X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"80",X"8A",X"80",
		X"B7",X"20",X"01",X"1C",X"AF",X"C6",X"28",X"EB",X"45",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",
		X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"80",X"B7",X"20",X"01",X"1C",X"AF",X"CB",
		X"08",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",
		X"A6",X"80",X"B7",X"20",X"01",X"1C",X"AF",X"C6",X"08",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",
		X"F7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"A6",X"45",X"8A",X"78",X"B7",X"20",X"01",X"1C",
		X"AF",X"39",X"8E",X"84",X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",X"B5",X"03",X"E3",X"26",X"03",
		X"7E",X"93",X"35",X"A6",X"44",X"2A",X"69",X"AE",X"48",X"EC",X"81",X"D7",X"00",X"AF",X"E3",X"8E",
		X"88",X"C8",X"48",X"AE",X"86",X"EC",X"81",X"97",X"01",X"D7",X"02",X"A6",X"84",X"43",X"97",X"04",
		X"C1",X"60",X"25",X"21",X"C1",X"78",X"22",X"1D",X"8E",X"01",X"20",X"A6",X"45",X"84",X"07",X"A6",
		X"86",X"84",X"07",X"9B",X"02",X"84",X"1F",X"8E",X"93",X"C2",X"A6",X"86",X"27",X"07",X"96",X"00",
		X"BB",X"03",X"EA",X"97",X"00",X"96",X"01",X"81",X"01",X"26",X"0A",X"A6",X"45",X"84",X"07",X"97",
		X"02",X"DB",X"02",X"D7",X"02",X"86",X"01",X"1F",X"01",X"96",X"00",X"E6",X"84",X"D4",X"04",X"E7",
		X"84",X"AA",X"84",X"A7",X"84",X"AE",X"E1",X"E6",X"80",X"E7",X"44",X"AF",X"48",X"1C",X"F3",X"39",
		X"AE",X"48",X"E6",X"02",X"C4",X"7F",X"E7",X"44",X"30",X"03",X"AF",X"48",X"30",X"1D",X"CC",X"00",
		X"00",X"DD",X"05",X"20",X"11",X"AE",X"48",X"E6",X"02",X"E7",X"44",X"30",X"03",X"AF",X"48",X"30",
		X"1D",X"CC",X"01",X"00",X"DD",X"05",X"EC",X"84",X"D7",X"00",X"8E",X"88",X"C8",X"48",X"AE",X"86",
		X"EC",X"81",X"97",X"01",X"D7",X"02",X"A6",X"84",X"43",X"97",X"04",X"96",X"05",X"27",X"25",X"C1",
		X"60",X"25",X"21",X"C1",X"78",X"22",X"1D",X"8E",X"01",X"20",X"A6",X"45",X"84",X"07",X"A6",X"86",
		X"84",X"07",X"9B",X"02",X"84",X"1F",X"8E",X"93",X"C2",X"A6",X"86",X"27",X"07",X"96",X"00",X"BB",
		X"03",X"EA",X"97",X"00",X"96",X"01",X"81",X"01",X"26",X"0A",X"A6",X"45",X"84",X"07",X"97",X"02",
		X"DB",X"02",X"D7",X"02",X"4F",X"1F",X"01",X"DC",X"05",X"27",X"02",X"30",X"8B",X"96",X"00",X"E6",
		X"84",X"D4",X"04",X"E7",X"84",X"AA",X"84",X"A7",X"84",X"1A",X"50",X"F6",X"20",X"01",X"2B",X"FB",
		X"D6",X"02",X"F7",X"20",X"00",X"F6",X"20",X"01",X"2B",X"FB",X"B7",X"20",X"01",X"1C",X"AF",X"1C",
		X"F3",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"8E",X"84",X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",X"B5",X"03",X"E3",X"26",X"03",
		X"7E",X"94",X"62",X"A6",X"44",X"2B",X"03",X"7E",X"94",X"4D",X"AE",X"48",X"EC",X"81",X"AF",X"E3",
		X"8E",X"88",X"C8",X"48",X"AE",X"86",X"EC",X"81",X"97",X"01",X"D7",X"02",X"A6",X"84",X"97",X"04",
		X"96",X"01",X"81",X"01",X"26",X"0A",X"A6",X"45",X"84",X"07",X"97",X"02",X"DB",X"02",X"D7",X"02",
		X"86",X"01",X"1F",X"01",X"E6",X"84",X"D4",X"04",X"DB",X"00",X"25",X"06",X"03",X"04",X"D5",X"04",
		X"27",X"06",X"03",X"04",X"DA",X"04",X"03",X"04",X"A6",X"84",X"94",X"04",X"A7",X"84",X"EA",X"84",
		X"E7",X"84",X"AE",X"E1",X"E6",X"80",X"E7",X"44",X"AF",X"48",X"1C",X"F3",X"39",X"AE",X"48",X"E6",
		X"02",X"C4",X"7F",X"E7",X"44",X"30",X"03",X"AF",X"48",X"30",X"1D",X"CC",X"00",X"00",X"DD",X"05",
		X"20",X"11",X"AE",X"48",X"E6",X"02",X"E7",X"44",X"30",X"03",X"AF",X"48",X"30",X"1D",X"CC",X"01",
		X"00",X"DD",X"05",X"EC",X"84",X"D7",X"00",X"8E",X"88",X"C8",X"48",X"AE",X"86",X"EC",X"81",X"97",
		X"01",X"D7",X"02",X"A6",X"84",X"97",X"04",X"96",X"01",X"81",X"01",X"26",X"0A",X"A6",X"45",X"84",
		X"07",X"97",X"02",X"DB",X"02",X"D7",X"02",X"4F",X"1F",X"01",X"DC",X"05",X"27",X"02",X"30",X"8B",
		X"E6",X"84",X"D4",X"04",X"DB",X"00",X"25",X"06",X"03",X"04",X"D5",X"04",X"27",X"06",X"03",X"04",
		X"DA",X"04",X"03",X"04",X"A6",X"84",X"94",X"04",X"A7",X"84",X"EA",X"84",X"E7",X"84",X"1A",X"50",
		X"B6",X"20",X"01",X"2B",X"FB",X"96",X"02",X"B7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"F7",
		X"20",X"01",X"1C",X"AF",X"1C",X"F3",X"39",X"8E",X"84",X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",
		X"B5",X"03",X"E3",X"26",X"03",X"7E",X"95",X"52",X"A6",X"44",X"2B",X"03",X"7E",X"95",X"3D",X"AE",
		X"48",X"EC",X"81",X"AF",X"E3",X"8E",X"88",X"C8",X"48",X"AE",X"86",X"EC",X"81",X"97",X"01",X"D7",
		X"02",X"A6",X"84",X"97",X"04",X"96",X"01",X"81",X"01",X"26",X"0A",X"A6",X"45",X"84",X"07",X"97",
		X"02",X"DB",X"02",X"D7",X"02",X"86",X"01",X"1F",X"01",X"E6",X"84",X"D4",X"04",X"D0",X"00",X"2B",
		X"06",X"03",X"04",X"D5",X"04",X"27",X"01",X"5F",X"A6",X"84",X"94",X"04",X"A7",X"84",X"EA",X"84",
		X"E7",X"84",X"AE",X"E1",X"E6",X"80",X"E7",X"44",X"AF",X"48",X"1C",X"F3",X"39",X"AE",X"48",X"E6",
		X"02",X"C4",X"7F",X"E7",X"44",X"30",X"03",X"AF",X"48",X"30",X"1D",X"CC",X"00",X"00",X"DD",X"05",
		X"20",X"11",X"AE",X"48",X"E6",X"02",X"E7",X"44",X"30",X"03",X"AF",X"48",X"30",X"1D",X"CC",X"01",
		X"00",X"DD",X"05",X"EC",X"84",X"D7",X"00",X"8E",X"88",X"C8",X"48",X"AE",X"86",X"EC",X"81",X"97",
		X"01",X"D7",X"02",X"A6",X"84",X"97",X"04",X"96",X"01",X"81",X"01",X"26",X"0A",X"A6",X"45",X"84",
		X"07",X"97",X"02",X"DB",X"02",X"D7",X"02",X"4F",X"1F",X"01",X"DC",X"05",X"27",X"02",X"30",X"8B",
		X"E6",X"84",X"D4",X"04",X"D0",X"00",X"2B",X"06",X"03",X"04",X"D5",X"04",X"27",X"01",X"5F",X"A6",
		X"84",X"94",X"04",X"A7",X"84",X"EA",X"84",X"E7",X"84",X"1A",X"50",X"B6",X"20",X"01",X"2B",X"FB",
		X"96",X"02",X"B7",X"20",X"00",X"B6",X"20",X"01",X"2B",X"FB",X"F7",X"20",X"01",X"1C",X"AF",X"1C",
		X"F3",X"39",X"AE",X"48",X"A6",X"C8",X"12",X"27",X"03",X"7E",X"96",X"5B",X"6C",X"C8",X"12",X"E6",
		X"84",X"58",X"AF",X"E3",X"8E",X"88",X"C8",X"AE",X"85",X"EC",X"81",X"81",X"01",X"26",X"0A",X"A6",
		X"45",X"84",X"07",X"B7",X"00",X"00",X"FB",X"00",X"00",X"E7",X"C8",X"10",X"A6",X"84",X"A7",X"C8",
		X"11",X"AE",X"E1",X"EC",X"02",X"ED",X"4E",X"A6",X"04",X"A7",X"4A",X"30",X"05",X"9F",X"07",X"9E",
		X"12",X"EC",X"84",X"DD",X"12",X"34",X"10",X"CC",X"00",X"13",X"BD",X"82",X"17",X"35",X"10",X"A6",
		X"45",X"97",X"0D",X"DF",X"09",X"EC",X"C4",X"DD",X"0B",X"AF",X"C4",X"1F",X"13",X"9E",X"09",X"A6",
		X"04",X"2A",X"08",X"9E",X"07",X"A6",X"80",X"A7",X"44",X"20",X"08",X"9E",X"07",X"A6",X"80",X"84",
		X"7F",X"A7",X"44",X"AF",X"48",X"96",X"0D",X"A7",X"45",X"34",X"40",X"DE",X"09",X"EC",X"46",X"AE",
		X"4C",X"35",X"40",X"ED",X"46",X"AF",X"4C",X"EF",X"E3",X"DE",X"0B",X"35",X"06",X"ED",X"42",X"1F",
		X"03",X"DC",X"0B",X"ED",X"C4",X"DC",X"09",X"ED",X"42",X"1F",X"03",X"8E",X"84",X"B9",X"A6",X"45",
		X"84",X"07",X"A6",X"86",X"B5",X"03",X"E3",X"26",X"03",X"7E",X"96",X"C5",X"AE",X"48",X"A6",X"44",
		X"2B",X"03",X"7E",X"97",X"2E",X"E6",X"01",X"2B",X"25",X"D7",X"00",X"86",X"01",X"E6",X"C8",X"10",
		X"1F",X"01",X"A6",X"84",X"A4",X"C8",X"11",X"9B",X"00",X"25",X"08",X"63",X"C8",X"11",X"A5",X"C8",
		X"11",X"27",X"24",X"63",X"C8",X"11",X"A4",X"C8",X"11",X"63",X"C8",X"11",X"20",X"19",X"D7",X"00",
		X"86",X"01",X"E6",X"C8",X"10",X"1F",X"01",X"A6",X"84",X"A4",X"C8",X"11",X"9B",X"00",X"63",X"C8",
		X"11",X"A5",X"C8",X"11",X"27",X"01",X"4F",X"E6",X"84",X"E4",X"C8",X"11",X"E7",X"84",X"AA",X"84",
		X"A7",X"84",X"7E",X"97",X"90",X"AE",X"48",X"E6",X"01",X"2B",X"25",X"D7",X"00",X"86",X"01",X"E6",
		X"C8",X"10",X"1F",X"01",X"A6",X"84",X"A4",X"C8",X"11",X"9B",X"00",X"25",X"08",X"63",X"C8",X"11",
		X"A5",X"C8",X"11",X"27",X"24",X"63",X"C8",X"11",X"A4",X"C8",X"11",X"63",X"C8",X"11",X"20",X"19",
		X"D7",X"00",X"86",X"01",X"E6",X"C8",X"10",X"1F",X"01",X"A6",X"84",X"A4",X"C8",X"11",X"9B",X"00",
		X"63",X"C8",X"11",X"A5",X"C8",X"11",X"27",X"01",X"4F",X"E6",X"84",X"E4",X"C8",X"11",X"E7",X"84",
		X"AA",X"84",X"A7",X"84",X"1A",X"50",X"F6",X"20",X"01",X"2B",X"FB",X"E6",X"C8",X"10",X"F7",X"20",
		X"00",X"F6",X"20",X"01",X"2B",X"FB",X"B7",X"20",X"01",X"1C",X"AF",X"7E",X"97",X"90",X"E6",X"01",
		X"2B",X"24",X"D7",X"00",X"4F",X"E6",X"C8",X"10",X"1F",X"01",X"A6",X"84",X"A4",X"C8",X"11",X"9B",
		X"00",X"25",X"08",X"63",X"C8",X"11",X"A5",X"C8",X"11",X"27",X"23",X"63",X"C8",X"11",X"A4",X"C8",
		X"11",X"63",X"C8",X"11",X"20",X"18",X"D7",X"00",X"4F",X"E6",X"C8",X"10",X"1F",X"01",X"A6",X"84",
		X"A4",X"C8",X"11",X"9B",X"00",X"63",X"C8",X"11",X"A5",X"C8",X"11",X"27",X"01",X"4F",X"E6",X"84",
		X"E4",X"C8",X"11",X"E7",X"84",X"AA",X"84",X"A7",X"84",X"1A",X"50",X"F6",X"20",X"01",X"2B",X"FB",
		X"E6",X"C8",X"10",X"F7",X"20",X"00",X"F6",X"20",X"01",X"2B",X"FB",X"B7",X"20",X"01",X"1C",X"AF",
		X"A6",X"4A",X"4A",X"26",X"09",X"6F",X"C8",X"12",X"BD",X"98",X"C2",X"86",X"80",X"39",X"A7",X"4A",
		X"EC",X"4E",X"E3",X"46",X"ED",X"46",X"63",X"C8",X"11",X"4F",X"39",X"96",X"20",X"2B",X"03",X"7E",
		X"97",X"EC",X"AE",X"48",X"A6",X"80",X"81",X"FF",X"26",X"0C",X"BD",X"98",X"C2",X"CC",X"00",X"00",
		X"FD",X"03",X"E7",X"1A",X"08",X"39",X"AF",X"48",X"8E",X"99",X"6D",X"48",X"AE",X"86",X"EC",X"02",
		X"DD",X"1D",X"A6",X"01",X"34",X"02",X"A6",X"84",X"8E",X"98",X"E4",X"30",X"86",X"A6",X"02",X"97",
		X"1F",X"10",X"AE",X"84",X"35",X"02",X"E6",X"A0",X"86",X"08",X"DD",X"20",X"CC",X"00",X"10",X"ED",
		X"46",X"1C",X"F7",X"1A",X"04",X"39",X"8E",X"84",X"B9",X"A6",X"45",X"84",X"07",X"A6",X"86",X"B5",
		X"03",X"E3",X"27",X"08",X"A6",X"44",X"2B",X"04",X"86",X"7F",X"20",X"02",X"86",X"FF",X"B7",X"00",
		X"00",X"AE",X"48",X"EC",X"46",X"E3",X"81",X"ED",X"46",X"A6",X"80",X"B4",X"00",X"00",X"A7",X"44",
		X"AF",X"48",X"4F",X"39",X"98",X"2C",X"98",X"32",X"98",X"38",X"98",X"3E",X"98",X"44",X"98",X"48",
		X"98",X"4C",X"98",X"44",X"98",X"48",X"98",X"4C",X"98",X"44",X"98",X"48",X"98",X"4C",X"98",X"44",
		X"98",X"48",X"98",X"4C",X"01",X"02",X"03",X"04",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",
		X"9E",X"12",X"34",X"10",X"30",X"02",X"CC",X"00",X"11",X"BD",X"82",X"17",X"35",X"10",X"EC",X"84",
		X"27",X"5F",X"DD",X"12",X"34",X"10",X"30",X"02",X"34",X"10",X"9E",X"10",X"30",X"02",X"34",X"10",
		X"EC",X"84",X"10",X"93",X"10",X"27",X"26",X"8E",X"03",X"F1",X"ED",X"84",X"35",X"06",X"ED",X"02",
		X"35",X"06",X"ED",X"04",X"35",X"06",X"ED",X"06",X"ED",X"94",X"ED",X"98",X"02",X"EC",X"84",X"ED",
		X"98",X"04",X"EC",X"02",X"83",X"00",X"02",X"ED",X"98",X"06",X"AE",X"06",X"39",X"8E",X"03",X"F1",
		X"ED",X"84",X"35",X"06",X"ED",X"02",X"35",X"06",X"ED",X"04",X"35",X"06",X"ED",X"06",X"ED",X"98",
		X"02",X"DD",X"0E",X"ED",X"98",X"04",X"EC",X"02",X"83",X"00",X"02",X"ED",X"98",X"06",X"AE",X"06",
		X"39",X"39",X"AE",X"C4",X"11",X"93",X"0E",X"26",X"0A",X"9F",X"0E",X"9C",X"10",X"26",X"0C",X"AF",
		X"02",X"20",X"08",X"EC",X"42",X"34",X"06",X"AF",X"F1",X"ED",X"02",X"DC",X"12",X"DF",X"12",X"ED",
		X"C4",X"1F",X"13",X"39",X"80",X"45",X"01",X"8F",X"DC",X"01",X"9C",X"8D",X"01",X"A7",X"8E",X"01",
		X"B8",X"8F",X"01",X"BD",X"90",X"01",X"C5",X"91",X"01",X"CE",X"F2",X"01",X"E4",X"33",X"01",X"F1",
		X"94",X"01",X"80",X"45",X"02",X"8C",X"44",X"02",X"91",X"85",X"02",X"AE",X"84",X"02",X"B4",X"35",
		X"02",X"BA",X"46",X"02",X"BF",X"77",X"02",X"CD",X"78",X"02",X"DE",X"79",X"02",X"99",X"45",X"99",
		X"47",X"99",X"49",X"99",X"4B",X"99",X"4D",X"99",X"4F",X"99",X"51",X"99",X"53",X"99",X"55",X"99",
		X"57",X"99",X"59",X"99",X"5B",X"99",X"5D",X"99",X"5F",X"99",X"61",X"99",X"63",X"99",X"65",X"99",
		X"67",X"99",X"69",X"99",X"6B",X"00",X"FF",X"01",X"FF",X"02",X"FF",X"03",X"FF",X"04",X"FF",X"05",
		X"FF",X"06",X"FF",X"07",X"FF",X"08",X"FF",X"09",X"FF",X"0A",X"FF",X"0B",X"FF",X"0A",X"FF",X"0D",
		X"FF",X"0E",X"FF",X"0F",X"FF",X"10",X"FF",X"11",X"FF",X"12",X"FF",X"13",X"FF",X"99",X"95",X"99",
		X"99",X"99",X"9D",X"99",X"A1",X"99",X"A5",X"99",X"A9",X"99",X"AD",X"99",X"B1",X"99",X"B5",X"99",
		X"B9",X"99",X"BD",X"99",X"C1",X"99",X"C5",X"99",X"C9",X"99",X"CD",X"99",X"D1",X"99",X"D5",X"99",
		X"D9",X"99",X"DD",X"99",X"E1",X"00",X"00",X"8F",X"DC",X"03",X"00",X"9C",X"8D",X"06",X"00",X"A7",
		X"8E",X"09",X"00",X"B8",X"8F",X"0C",X"00",X"BD",X"90",X"0F",X"00",X"C5",X"91",X"12",X"00",X"CE",
		X"F2",X"15",X"00",X"E4",X"33",X"18",X"00",X"F1",X"94",X"1B",X"00",X"F9",X"25",X"1E",X"00",X"8C",
		X"44",X"21",X"00",X"91",X"85",X"1E",X"00",X"8C",X"44",X"24",X"00",X"AE",X"84",X"27",X"00",X"B4",
		X"35",X"2A",X"00",X"BA",X"46",X"2D",X"00",X"BF",X"77",X"30",X"00",X"CD",X"78",X"33",X"00",X"DE",
		X"79",X"36",X"00",X"F2",X"7A",X"E9",X"50",X"3A",X"68",X"3C",X"35",X"0D",X"0A",X"10",X"00",X"1F",
		X"59",X"95",X"9F",X"94",X"96",X"9C",X"8E",X"C0",X"40",X"C6",X"84",X"07",X"4F",X"47",X"23",X"E9",
		X"50",X"3A",X"68",X"3C",X"35",X"0D",X"0A",X"10",X"00",X"1F",X"59",X"95",X"9F",X"94",X"96",X"9C",
		X"8E",X"C0",X"40",X"C6",X"88",X"07",X"4F",X"47",X"23",X"E9",X"50",X"3A",X"68",X"3C",X"35",X"0D",
		X"0A",X"10",X"00",X"1F",X"59",X"95",X"9F",X"94",X"96",X"9C",X"8E",X"C0",X"40",X"C6",X"8A",X"07",
		X"4F",X"47",X"23",X"C0",X"50",X"31",X"31",X"61",X"31",X"1F",X"18",X"14",X"00",X"5F",X"1C",X"5F",
		X"5F",X"06",X"06",X"06",X"12",X"00",X"00",X"00",X"08",X"F6",X"F8",X"F9",X"08",X"ED",X"60",X"65",
		X"61",X"36",X"00",X"13",X"05",X"28",X"00",X"1F",X"02",X"1F",X"02",X"13",X"0C",X"19",X"1F",X"07",
		X"00",X"00",X"00",X"F6",X"04",X"E4",X"04",X"E9",X"10",X"62",X"60",X"01",X"60",X"11",X"15",X"15",
		X"00",X"11",X"12",X"11",X"16",X"0A",X"06",X"1F",X"1F",X"C2",X"02",X"00",X"80",X"31",X"81",X"01",
		X"04",X"E0",X"60",X"31",X"31",X"31",X"31",X"23",X"18",X"18",X"00",X"1F",X"1F",X"1F",X"1F",X"06",
		X"1F",X"1F",X"1F",X"02",X"02",X"02",X"02",X"FF",X"0F",X"0F",X"0F",X"E5",X"62",X"10",X"22",X"42",
		X"32",X"11",X"00",X"00",X"00",X"1D",X"3F",X"5F",X"1F",X"10",X"06",X"09",X"03",X"0F",X"0F",X"0F",
		X"0F",X"F7",X"57",X"37",X"F7",X"FC",X"60",X"35",X"3A",X"31",X"31",X"22",X"2C",X"00",X"00",X"56",
		X"5C",X"5C",X"5C",X"0E",X"11",X"11",X"11",X"09",X"06",X"0A",X"0A",X"46",X"36",X"35",X"35",X"FA",
		X"60",X"05",X"04",X"62",X"62",X"1C",X"15",X"12",X"00",X"9F",X"5F",X"06",X"1B",X"88",X"8B",X"8A",
		X"8A",X"06",X"04",X"02",X"03",X"57",X"03",X"01",X"28",X"C8",X"50",X"63",X"31",X"31",X"31",X"28",
		X"24",X"14",X"00",X"10",X"1A",X"13",X"1B",X"0F",X"1F",X"1F",X"1F",X"05",X"07",X"08",X"03",X"33",
		X"03",X"05",X"0B",X"D4",X"00",X"11",X"71",X"31",X"31",X"15",X"14",X"00",X"00",X"1B",X"9F",X"1D",
		X"1D",X"08",X"0B",X"03",X"01",X"00",X"00",X"00",X"00",X"F7",X"47",X"17",X"17",X"ED",X"60",X"65",
		X"61",X"36",X"01",X"13",X"0F",X"28",X"09",X"1F",X"0A",X"1F",X"0A",X"13",X"0C",X"19",X"1F",X"07",
		X"08",X"09",X"0C",X"F6",X"04",X"E4",X"04",X"CA",X"60",X"3A",X"38",X"34",X"34",X"30",X"19",X"2D",
		X"00",X"09",X"1C",X"1F",X"1B",X"94",X"96",X"97",X"8D",X"12",X"10",X"0D",X"0C",X"57",X"03",X"01",
		X"08",X"C2",X"60",X"0A",X"08",X"68",X"68",X"32",X"2A",X"26",X"00",X"92",X"52",X"06",X"1F",X"88",
		X"8B",X"94",X"94",X"12",X"50",X"8D",X"CC",X"57",X"03",X"01",X"28",X"FD",X"FF",X"00",X"01",X"01",
		X"02",X"13",X"00",X"00",X"00",X"18",X"1B",X"1C",X"1A",X"14",X"14",X"13",X"12",X"19",X"93",X"82",
		X"D1",X"00",X"3B",X"3D",X"3F",X"FB",X"00",X"70",X"04",X"02",X"42",X"00",X"00",X"00",X"00",X"1F",
		X"1F",X"1F",X"1F",X"10",X"10",X"12",X"13",X"80",X"40",X"C0",X"80",X"DF",X"FF",X"FF",X"FF",X"EC",
		X"60",X"62",X"05",X"10",X"50",X"1A",X"16",X"00",X"00",X"1F",X"9F",X"1F",X"1F",X"16",X"13",X"1F",
		X"1F",X"80",X"D0",X"54",X"98",X"A9",X"A5",X"07",X"07",X"FD",X"00",X"01",X"01",X"01",X"01",X"12",
		X"00",X"00",X"00",X"1A",X"1A",X"1A",X"1A",X"0F",X"14",X"12",X"11",X"19",X"90",X"9D",X"FD",X"00",
		X"04",X"DD",X"FF",X"FB",X"00",X"4F",X"00",X"00",X"40",X"0B",X"00",X"00",X"06",X"1B",X"1B",X"1B",
		X"1B",X"14",X"14",X"15",X"17",X"80",X"40",X"C0",X"80",X"1F",X"FF",X"FF",X"FF",X"D0",X"50",X"63",
		X"31",X"31",X"31",X"1A",X"1A",X"1B",X"00",X"10",X"1A",X"13",X"1B",X"0F",X"1F",X"1F",X"1F",X"00",
		X"00",X"00",X"00",X"33",X"03",X"05",X"0B",X"C8",X"00",X"68",X"32",X"32",X"32",X"24",X"18",X"1F",
		X"00",X"10",X"1C",X"14",X"1F",X"0A",X"18",X"12",X"1A",X"0C",X"0A",X"02",X"01",X"33",X"03",X"05",
		X"0B",X"C8",X"50",X"68",X"34",X"32",X"32",X"22",X"20",X"1B",X"00",X"10",X"16",X"10",X"1F",X"0F",
		X"13",X"0A",X"1F",X"0C",X"0A",X"06",X"01",X"33",X"03",X"05",X"0B",X"D4",X"00",X"11",X"51",X"31",
		X"31",X"14",X"10",X"00",X"00",X"1B",X"14",X"1B",X"1B",X"0C",X"0A",X"13",X"11",X"00",X"00",X"00",
		X"00",X"F7",X"F7",X"17",X"17",X"ED",X"60",X"65",X"61",X"36",X"00",X"13",X"05",X"28",X"00",X"1F",
		X"12",X"13",X"14",X"13",X"0C",X"19",X"1F",X"07",X"00",X"00",X"00",X"F6",X"04",X"E4",X"04",X"E2",
		X"10",X"6B",X"67",X"03",X"62",X"0C",X"0A",X"08",X"00",X"12",X"18",X"0F",X"11",X"0A",X"06",X"14",
		X"1F",X"00",X"00",X"00",X"00",X"21",X"51",X"01",X"06",X"E9",X"10",X"62",X"60",X"01",X"60",X"11",
		X"15",X"15",X"00",X"11",X"12",X"11",X"0C",X"0A",X"06",X"1F",X"1F",X"C2",X"02",X"00",X"91",X"31",
		X"81",X"01",X"F7",X"FD",X"00",X"71",X"40",X"01",X"01",X"1B",X"00",X"00",X"00",X"1F",X"14",X"13",
		X"14",X"00",X"0E",X"0F",X"0E",X"12",X"74",X"9D",X"19",X"0E",X"08",X"DD",X"FF",X"FD",X"00",X"71",
		X"40",X"01",X"01",X"06",X"00",X"00",X"00",X"1F",X"14",X"13",X"14",X"00",X"10",X"12",X"10",X"D2",
		X"74",X"9D",X"19",X"0E",X"08",X"DD",X"FF",X"FD",X"00",X"71",X"40",X"01",X"01",X"02",X"00",X"00",
		X"00",X"1F",X"0A",X"08",X"07",X"00",X"10",X"12",X"10",X"D2",X"74",X"9D",X"19",X"0E",X"08",X"DD",
		X"FF",X"C3",X"00",X"53",X"46",X"03",X"41",X"26",X"0C",X"1A",X"00",X"0F",X"1F",X"1F",X"1F",X"00",
		X"12",X"0B",X"0F",X"12",X"D4",X"9D",X"19",X"0E",X"08",X"DD",X"FF",X"C3",X"00",X"53",X"46",X"03",
		X"41",X"26",X"10",X"13",X"00",X"0F",X"1F",X"1F",X"1F",X"00",X"10",X"0B",X"0F",X"52",X"D4",X"9D",
		X"19",X"0E",X"08",X"DD",X"FF",X"C3",X"00",X"79",X"64",X"75",X"34",X"34",X"14",X"24",X"00",X"1F",
		X"0C",X"1F",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"7F",X"7F",X"7F",X"DD",
		X"FF",X"80",X"02",X"F1",X"13",X"00",X"00",X"00",X"00",X"0A",X"1F",X"1F",X"1F",X"00",X"00",X"0B",
		X"00",X"12",X"64",X"9D",X"19",X"0E",X"08",X"DD",X"FF",X"FE",X"FF",X"74",X"41",X"02",X"02",X"06",
		X"09",X"00",X"00",X"1F",X"0C",X"1F",X"1F",X"00",X"00",X"0B",X"00",X"12",X"64",X"9D",X"19",X"0E",
		X"08",X"DD",X"FF",X"E0",X"60",X"3A",X"32",X"35",X"31",X"16",X"17",X"20",X"00",X"1F",X"1F",X"15",
		X"1F",X"06",X"1F",X"1F",X"1F",X"02",X"02",X"02",X"02",X"FF",X"0F",X"0F",X"0F",X"FD",X"60",X"32",
		X"62",X"32",X"62",X"1D",X"1B",X"04",X"04",X"10",X"11",X"13",X"12",X"1F",X"1F",X"1F",X"1F",X"0B",
		X"00",X"00",X"00",X"07",X"08",X"09",X"08",X"FB",X"50",X"36",X"34",X"34",X"32",X"1D",X"27",X"2A",
		X"00",X"1F",X"1F",X"98",X"9F",X"0D",X"0E",X"0E",X"91",X"06",X"08",X"05",X"05",X"54",X"66",X"44",
		X"04",X"FA",X"60",X"02",X"62",X"12",X"32",X"1C",X"1F",X"24",X"08",X"9F",X"5B",X"90",X"50",X"09",
		X"1F",X"09",X"03",X"00",X"00",X"00",X"00",X"13",X"06",X"F5",X"06",X"FA",X"53",X"08",X"04",X"64",
		X"62",X"20",X"21",X"12",X"00",X"5B",X"1F",X"19",X"52",X"12",X"94",X"14",X"13",X"00",X"00",X"00",
		X"00",X"29",X"65",X"16",X"08",X"89",X"00",X"9D",X"F9",X"81",X"00",X"F0",X"88",X"9B",X"85",X"80",
		X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"21",
		X"00",X"00",X"78",X"00",X"81",X"00",X"F0",X"81",X"01",X"E0",X"88",X"9B",X"85",X"80",X"21",X"00",
		X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9B",X"85",X"80",X"2A",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"81",X"00",X"F0",X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",
		X"F0",X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"81",X"03",X"C0",
		X"81",X"00",X"F0",X"88",X"9B",X"85",X"80",X"2A",X"00",X"00",X"78",X"00",X"81",X"01",X"68",X"80",
		X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"81",X"00",X"78",X"88",X"9B",X"85",X"80",X"21",
		X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"78",X"00",
		X"81",X"00",X"F0",X"80",X"2E",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"81",X"02",X"D0",X"88",
		X"9B",X"85",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"81",X"03",X"C0",X"81",X"00",
		X"78",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"F0",X"88",X"9B",X"85",X"80",X"21",X"00",
		X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9B",X"85",X"80",X"2E",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"81",X"00",X"78",X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"01",
		X"E0",X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"81",X"00",X"78",
		X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"01",X"68",X"88",X"9B",X"85",X"80",
		X"2E",X"00",X"00",X"78",X"00",X"81",X"00",X"F0",X"81",X"00",X"78",X"88",X"9B",X"85",X"80",X"21",
		X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9B",X"85",X"80",X"1E",X"00",X"00",X"3C",X"00",
		X"80",X"1A",X"00",X"00",X"3C",X"00",X"81",X"01",X"E0",X"81",X"02",X"D0",X"80",X"21",X"00",X"00",
		X"78",X"00",X"81",X"03",X"48",X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",
		X"78",X"89",X"04",X"9F",X"35",X"81",X"00",X"50",X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"50",
		X"00",X"81",X"00",X"50",X"8A",X"81",X"01",X"E0",X"80",X"21",X"00",X"00",X"3C",X"00",X"80",X"21",
		X"00",X"00",X"3C",X"00",X"80",X"1E",X"00",X"00",X"3C",X"00",X"80",X"1E",X"00",X"00",X"3C",X"00",
		X"80",X"1A",X"00",X"00",X"3C",X"00",X"80",X"1A",X"00",X"00",X"3C",X"00",X"80",X"18",X"00",X"00",
		X"3C",X"00",X"80",X"18",X"00",X"00",X"3C",X"00",X"8A",X"89",X"00",X"9F",X"7D",X"88",X"9A",X"9B",
		X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",
		X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",
		X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"99",X"FF",X"80",X"58",X"00",X"00",
		X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"21",
		X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",
		X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",
		X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",
		X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",X"00",
		X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"10",X"80",X"21",X"00",X"00",
		X"F0",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",
		X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"99",X"FF",X"80",X"6C",X"00",
		X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",
		X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",
		X"08",X"97",X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",
		X"94",X"12",X"2A",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"2A",X"00",X"00",X"78",X"00",X"88",
		X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",
		X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"0F",X"10",X"80",X"21",X"00",X"00",X"F0",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",
		X"12",X"FF",X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",
		X"30",X"97",X"12",X"FF",X"00",X"0F",X"08",X"97",X"12",X"FF",X"00",X"50",X"03",X"80",X"30",X"00",
		X"00",X"F0",X"00",X"88",X"99",X"FF",X"80",X"6C",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",
		X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9A",
		X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",
		X"81",X"00",X"F0",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"10",X"80",
		X"21",X"00",X"00",X"F0",X"00",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"07",X"10",X"80",X"21",
		X"00",X"00",X"78",X"00",X"88",X"99",X"E5",X"80",X"6C",X"00",X"01",X"68",X"00",X"88",X"9A",X"9B",
		X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",
		X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",
		X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",
		X"12",X"FF",X"00",X"0F",X"10",X"80",X"21",X"00",X"00",X"F0",X"00",X"88",X"99",X"FF",X"80",X"6C",
		X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",
		X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",
		X"07",X"08",X"97",X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9A",
		X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",
		X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"21",X"00",X"00",
		X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",
		X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",
		X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",
		X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",
		X"00",X"88",X"9B",X"6B",X"94",X"12",X"2E",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"2E",X"00",
		X"00",X"78",X"00",X"88",X"99",X"FF",X"80",X"5A",X"00",X"00",X"78",X"00",X"88",X"9A",X"9B",X"94",
		X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"10",X"80",X"21",X"00",X"00",X"F0",X"00",X"88",X"9B",
		X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",X"03",
		X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",
		X"0F",X"10",X"80",X"21",X"00",X"00",X"F0",X"00",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"07",
		X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"99",X"FF",X"80",X"5A",X"00",X"00",
		X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"19",X"80",X"5C",X"00",X"00",X"3C",X"00",X"80",X"5C",
		X"00",X"00",X"3C",X"00",X"80",X"5C",X"00",X"00",X"78",X"00",X"88",X"99",X"E5",X"80",X"6C",X"00",
		X"02",X"58",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"07",X"10",X"80",
		X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",
		X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",
		X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",
		X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"21",X"00",
		X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",
		X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",
		X"2E",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"2E",X"00",X"00",X"78",X"00",X"88",X"99",X"FF",
		X"80",X"5A",X"00",X"00",X"78",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",
		X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",
		X"FF",X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",
		X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",
		X"78",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"10",X"80",X"21",
		X"00",X"00",X"F0",X"00",X"88",X"99",X"FF",X"80",X"6C",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",
		X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",
		X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",
		X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",
		X"12",X"FF",X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",
		X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",
		X"00",X"78",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"10",X"80",
		X"21",X"00",X"00",X"F0",X"00",X"88",X"9B",X"6B",X"94",X"12",X"2E",X"97",X"12",X"FF",X"00",X"0F",
		X"08",X"80",X"2E",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",
		X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",
		X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",
		X"00",X"81",X"00",X"78",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",
		X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",
		X"07",X"08",X"97",X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"94",X"12",
		X"1E",X"97",X"12",X"FF",X"00",X"07",X"08",X"80",X"1E",X"00",X"00",X"3C",X"00",X"94",X"12",X"1A",
		X"97",X"12",X"FF",X"00",X"07",X"08",X"80",X"1A",X"00",X"00",X"3C",X"00",X"88",X"9A",X"9B",X"94",
		X"12",X"21",X"97",X"12",X"FF",X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"99",
		X"E5",X"80",X"6C",X"00",X"01",X"68",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"99",X"FF",X"89",X"05",X"A4",X"D0",
		X"80",X"6C",X"00",X"00",X"78",X"00",X"8A",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"0F",X"08",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"99",X"E5",X"80",X"5C",X"00",X"01",
		X"E0",X"00",X"88",X"9A",X"19",X"80",X"6C",X"00",X"00",X"F0",X"00",X"80",X"6C",X"00",X"00",X"78",
		X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0F",X"08",X"80",X"21",X"00",
		X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",
		X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9B",X"B9",X"94",X"12",
		X"30",X"97",X"12",X"FF",X"00",X"00",X"08",X"97",X"12",X"FF",X"00",X"1A",X"03",X"80",X"30",X"00",
		X"00",X"50",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",X"0A",X"08",X"80",
		X"21",X"00",X"00",X"50",X"00",X"88",X"99",X"FF",X"80",X"6C",X"00",X"00",X"50",X"00",X"88",X"9B",
		X"B9",X"94",X"12",X"2E",X"97",X"12",X"FF",X"00",X"00",X"08",X"97",X"12",X"FF",X"00",X"1A",X"03",
		X"80",X"2E",X"00",X"00",X"50",X"00",X"88",X"9B",X"6B",X"94",X"12",X"2E",X"97",X"12",X"FF",X"00",
		X"0A",X"08",X"80",X"2E",X"00",X"00",X"50",X"00",X"88",X"99",X"FF",X"80",X"65",X"00",X"00",X"50",
		X"00",X"88",X"9B",X"B9",X"94",X"12",X"2D",X"97",X"12",X"FF",X"00",X"00",X"08",X"97",X"12",X"FF",
		X"00",X"1A",X"03",X"80",X"2D",X"00",X"00",X"50",X"00",X"88",X"9B",X"6B",X"94",X"12",X"2A",X"97",
		X"12",X"FF",X"00",X"0A",X"08",X"80",X"2A",X"00",X"00",X"50",X"00",X"88",X"99",X"FF",X"80",X"61",
		X"00",X"00",X"50",X"00",X"88",X"9B",X"B9",X"94",X"12",X"2C",X"97",X"12",X"FF",X"00",X"00",X"08",
		X"97",X"12",X"FF",X"00",X"1A",X"03",X"80",X"2C",X"00",X"00",X"50",X"00",X"88",X"9B",X"6B",X"94",
		X"12",X"28",X"97",X"12",X"FF",X"00",X"0A",X"08",X"80",X"28",X"00",X"00",X"50",X"00",X"88",X"99",
		X"FF",X"80",X"5C",X"00",X"00",X"50",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"07",X"10",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"99",X"FF",X"89",X"06",X"A6",X"10",
		X"80",X"6C",X"00",X"00",X"3C",X"00",X"8A",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"07",X"08",X"80",X"21",X"00",X"00",X"3C",X"00",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",
		X"07",X"08",X"80",X"21",X"00",X"00",X"3C",X"00",X"94",X"12",X"1E",X"97",X"12",X"FF",X"00",X"07",
		X"08",X"80",X"1E",X"00",X"00",X"3C",X"00",X"94",X"12",X"1E",X"97",X"12",X"FF",X"00",X"07",X"08",
		X"80",X"1E",X"00",X"00",X"3C",X"00",X"94",X"12",X"1A",X"97",X"12",X"FF",X"00",X"07",X"08",X"80",
		X"1A",X"00",X"00",X"3C",X"00",X"94",X"12",X"1A",X"97",X"12",X"FF",X"00",X"07",X"08",X"80",X"1A",
		X"00",X"00",X"3C",X"00",X"94",X"12",X"18",X"97",X"12",X"FF",X"00",X"07",X"08",X"80",X"18",X"00",
		X"00",X"3C",X"00",X"94",X"12",X"18",X"97",X"12",X"FF",X"00",X"07",X"08",X"80",X"18",X"00",X"00",
		X"3C",X"00",X"8A",X"88",X"9A",X"B5",X"89",X"00",X"A6",X"9A",X"89",X"03",X"A6",X"9E",X"80",X"2A",
		X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",
		X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",
		X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"8A",X"81",
		X"00",X"78",X"80",X"3D",X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",X"00",X"80",X"3D",
		X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",
		X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",
		X"3C",X"00",X"80",X"34",X"00",X"00",X"3C",X"00",X"89",X"03",X"A7",X"0C",X"80",X"3A",X"00",X"00",
		X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3A",
		X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",
		X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"8A",X"81",X"00",X"78",
		X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"28",
		X"00",X"00",X"3C",X"00",X"80",X"2A",X"00",X"00",X"3C",X"00",X"80",X"2C",X"00",X"00",X"3C",X"00",
		X"80",X"2E",X"00",X"00",X"3C",X"00",X"89",X"03",X"A7",X"7A",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",
		X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"36",X"00",X"00",X"78",X"00",X"80",X"31",
		X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"8A",X"81",X"00",X"F0",X"89",X"02",
		X"A7",X"B2",X"80",X"32",X"00",X"00",X"3C",X"00",X"80",X"34",X"00",X"00",X"3C",X"00",X"80",X"38",
		X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"00",X"3C",X"00",X"80",X"3D",X"00",X"00",X"3C",X"00",
		X"80",X"3E",X"00",X"00",X"3C",X"00",X"8A",X"89",X"03",X"A7",X"DB",X"80",X"2A",X"00",X"00",X"78",
		X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"34",X"00",
		X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",
		X"31",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"8A",X"80",X"40",X"00",X"00",
		X"3C",X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",X"80",X"48",X"00",X"00",X"3C",X"00",X"80",X"3A",
		X"00",X"00",X"3C",X"00",X"80",X"48",X"00",X"00",X"3C",X"00",X"80",X"46",X"00",X"00",X"3C",X"00",
		X"80",X"41",X"00",X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",X"80",X"48",X"00",X"00",
		X"3C",X"00",X"80",X"3A",X"00",X"00",X"3C",X"00",X"80",X"42",X"00",X"00",X"3C",X"00",X"80",X"44",
		X"00",X"00",X"3C",X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"3C",X"00",
		X"80",X"3E",X"00",X"00",X"3C",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",
		X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"31",
		X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"29",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",
		X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"38",
		X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",
		X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",
		X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"39",X"00",X"00",X"78",X"00",X"80",X"38",
		X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",
		X"80",X"31",X"00",X"00",X"78",X"00",X"81",X"00",X"F0",X"80",X"45",X"00",X"00",X"3C",X"00",X"80",
		X"41",X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"00",X"3C",
		X"00",X"80",X"31",X"00",X"00",X"F0",X"00",X"81",X"00",X"F0",X"80",X"25",X"00",X"00",X"78",X"00",
		X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",
		X"00",X"00",X"78",X"00",X"80",X"29",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",
		X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",
		X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"35",
		X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"39",X"00",X"00",
		X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"2E",
		X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"89",X"03",X"A9",X"AE",X"81",X"00",
		X"78",X"80",X"2E",X"00",X"00",X"3C",X"00",X"80",X"31",X"00",X"00",X"3C",X"00",X"8A",X"80",X"35",
		X"00",X"00",X"3C",X"00",X"80",X"31",X"00",X"00",X"3C",X"00",X"80",X"2E",X"00",X"00",X"3C",X"00",
		X"80",X"2A",X"00",X"00",X"3C",X"00",X"89",X"03",X"A9",X"DA",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",
		X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3E",
		X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"8A",X"81",X"00",X"78",X"80",X"3D",
		X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",X"00",X"80",X"3D",X"00",X"00",X"78",X"00",
		X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",
		X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"3C",X"00",X"80",X"34",
		X"00",X"00",X"3C",X"00",X"89",X"03",X"AA",X"48",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"2A",
		X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",
		X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",
		X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"8A",X"81",X"00",X"78",X"80",X"3A",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"31",
		X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"3C",X"00",
		X"80",X"2A",X"00",X"00",X"3C",X"00",X"80",X"2C",X"00",X"00",X"3C",X"00",X"80",X"2E",X"00",X"00",
		X"3C",X"00",X"89",X"02",X"AA",X"B6",X"80",X"25",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",
		X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"38",
		X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"8A",X"80",X"25",X"00",X"00",X"78",
		X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",
		X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",
		X"3A",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",
		X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"24",X"00",
		X"00",X"78",X"00",X"81",X"00",X"F0",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",
		X"3C",X"00",X"80",X"2A",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"81",X"01",
		X"68",X"89",X"02",X"AB",X"45",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"36",X"00",X"00",X"78",X"00",X"80",X"32",X"00",
		X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"8A",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"36",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",
		X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",
		X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",
		X"78",X"00",X"81",X"00",X"F0",X"80",X"3D",X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",
		X"00",X"80",X"41",X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",X"00",X"80",X"3D",X"00",
		X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",X"00",X"80",X"48",X"00",X"00",X"3C",X"00",X"80",
		X"3E",X"00",X"00",X"3C",X"00",X"80",X"3D",X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",
		X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",X"00",X"89",X"03",X"AC",
		X"01",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",
		X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",
		X"36",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",
		X"00",X"8A",X"81",X"00",X"F0",X"89",X"02",X"AC",X"39",X"80",X"32",X"00",X"00",X"3C",X"00",X"80",
		X"34",X"00",X"00",X"3C",X"00",X"80",X"38",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"00",X"3C",
		X"00",X"80",X"3D",X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",X"00",X"8A",X"80",X"2A",
		X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",
		X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3D",X"00",X"00",
		X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"44",
		X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",X"00",
		X"80",X"48",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"48",X"00",X"00",
		X"78",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",X"44",
		X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",
		X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",
		X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"3D",
		X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",
		X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"3C",X"00",X"80",X"34",X"00",X"00",
		X"3C",X"00",X"80",X"42",X"00",X"00",X"3C",X"00",X"80",X"41",X"00",X"00",X"3C",X"00",X"80",X"3E",
		X"00",X"00",X"3C",X"00",X"80",X"38",X"00",X"00",X"3C",X"00",X"80",X"34",X"00",X"00",X"3C",X"00",
		X"80",X"32",X"00",X"00",X"3C",X"00",X"80",X"31",X"00",X"00",X"3C",X"00",X"80",X"2E",X"00",X"00",
		X"3C",X"00",X"90",X"8A",X"A6",X"93",X"9D",X"F5",X"B2",X"39",X"B6",X"B9",X"BB",X"63",X"AD",X"54",
		X"BB",X"74",X"9F",X"79",X"88",X"9A",X"33",X"89",X"04",X"AD",X"5B",X"81",X"2D",X"00",X"8A",X"89",
		X"00",X"AD",X"63",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",
		X"32",X"00",X"07",X"08",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",
		X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",
		X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"81",
		X"03",X"C0",X"80",X"36",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"36",
		X"00",X"02",X"58",X"00",X"80",X"38",X"00",X"00",X"F0",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",
		X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",
		X"78",X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"2C",
		X"00",X"03",X"48",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"81",X"03",X"C0",X"80",X"2A",X"00",X"00",X"F0",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",
		X"32",X"00",X"00",X"F0",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"F0",
		X"00",X"80",X"2A",X"00",X"00",X"F0",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"38",X"00",
		X"00",X"F0",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",
		X"2A",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",
		X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"3D",X"00",X"00",X"F0",X"00",X"80",X"3E",X"00",
		X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",
		X"38",X"00",X"00",X"F0",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",
		X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"42",X"00",X"00",X"F0",X"00",X"80",X"46",X"00",
		X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",
		X"48",X"00",X"00",X"78",X"00",X"80",X"46",X"00",X"00",X"F0",X"00",X"80",X"48",X"00",X"00",X"78",
		X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",
		X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"46",X"00",X"00",X"78",X"00",X"80",
		X"42",X"00",X"00",X"F0",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",
		X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",
		X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"F0",X"00",X"80",
		X"3E",X"00",X"00",X"78",X"00",X"80",X"40",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",
		X"00",X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"50",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",
		X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",
		X"4A",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"4D",X"00",X"00",X"3C",
		X"00",X"80",X"4E",X"00",X"00",X"3C",X"00",X"80",X"4E",X"00",X"07",X"F8",X"00",X"80",X"54",X"00",
		X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",X"80",X"45",X"00",X"00",X"78",X"00",X"80",
		X"49",X"00",X"00",X"78",X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",
		X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",X"4A",X"00",X"03",X"48",X"00",
		X"80",X"51",X"00",X"03",X"C0",X"00",X"80",X"4E",X"00",X"02",X"D0",X"00",X"80",X"55",X"00",X"00",
		X"78",X"00",X"80",X"49",X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"81",X"03",
		X"C0",X"80",X"38",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"06",X"CC",X"00",X"80",X"48",X"00",
		X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",X"80",X"54",X"00",X"01",X"68",X"00",X"80",
		X"4E",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"78",
		X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"04",X"38",X"00",X"80",X"4A",X"00",
		X"00",X"78",X"00",X"89",X"04",X"AF",X"D7",X"80",X"48",X"00",X"00",X"3C",X"00",X"80",X"4A",X"00",
		X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"8A",X"80",X"38",X"00",X"00",X"3C",X"00",
		X"80",X"3A",X"00",X"03",X"0C",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"89",X"04",X"B0",X"00",
		X"80",X"4D",X"00",X"00",X"3C",X"00",X"80",X"4E",X"00",X"00",X"3C",X"00",X"80",X"4E",X"00",X"00",
		X"78",X"00",X"8A",X"80",X"38",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"03",X"0C",X"00",X"81",
		X"00",X"78",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"4A",
		X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"78",X"00",
		X"80",X"4D",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"F0",X"00",X"80",X"48",X"00",X"00",
		X"3C",X"00",X"80",X"4A",X"00",X"03",X"0C",X"00",X"81",X"00",X"78",X"80",X"4A",X"00",X"00",X"78",
		X"00",X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"52",X"00",X"00",X"78",X"00",X"80",X"51",X"00",
		X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",
		X"4A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"81",X"00",X"78",X"80",X"4A",X"00",X"00",X"78",
		X"00",X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"4D",X"00",
		X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",
		X"4A",X"00",X"00",X"F0",X"00",X"80",X"3D",X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"03",X"0C",
		X"00",X"81",X"00",X"78",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",
		X"80",X"42",X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",
		X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"F0",X"00",X"80",X"4A",
		X"00",X"00",X"F0",X"00",X"80",X"51",X"00",X"00",X"F0",X"00",X"80",X"4E",X"00",X"00",X"F0",X"00",
		X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"52",X"00",X"00",X"78",X"00",X"80",X"54",X"00",X"00",
		X"78",X"00",X"80",X"52",X"00",X"07",X"08",X"00",X"80",X"54",X"00",X"00",X"78",X"00",X"80",X"48",
		X"00",X"00",X"78",X"00",X"80",X"52",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",
		X"80",X"45",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",
		X"78",X"00",X"81",X"03",X"C0",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",
		X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"F0",X"00",X"80",X"48",X"00",
		X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"F0",X"00",X"80",
		X"4A",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"F0",
		X"00",X"80",X"51",X"00",X"00",X"3C",X"00",X"80",X"52",X"00",X"00",X"3C",X"00",X"80",X"51",X"00",
		X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"3C",X"00",X"80",
		X"4E",X"00",X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",X"80",X"48",X"00",X"00",X"3C",
		X"00",X"80",X"4E",X"00",X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",X"80",X"48",X"00",
		X"00",X"3C",X"00",X"80",X"44",X"00",X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",X"80",
		X"44",X"00",X"00",X"3C",X"00",X"80",X"42",X"00",X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",X"3C",
		X"00",X"80",X"41",X"00",X"00",X"3C",X"00",X"80",X"4E",X"00",X"00",X"3C",X"00",X"80",X"44",X"00",
		X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"41",X"00",X"00",X"3C",X"00",X"80",X"44",X"00",X"00",
		X"3C",X"00",X"81",X"00",X"78",X"80",X"38",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"00",X"3C",
		X"00",X"81",X"00",X"78",X"80",X"4E",X"00",X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",
		X"80",X"44",X"00",X"00",X"3C",X"00",X"80",X"3E",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"00",
		X"3C",X"00",X"80",X"2A",X"00",X"00",X"3C",X"00",X"8A",X"88",X"9A",X"CF",X"89",X"00",X"B2",X"40",
		X"89",X"03",X"B2",X"44",X"81",X"01",X"E0",X"80",X"34",X"00",X"03",X"C0",X"00",X"80",X"3E",X"00",
		X"03",X"48",X"00",X"80",X"42",X"00",X"00",X"F0",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",
		X"38",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"8A",X"80",
		X"54",X"00",X"03",X"C0",X"00",X"80",X"48",X"00",X"04",X"B0",X"00",X"80",X"46",X"00",X"00",X"F0",
		X"00",X"80",X"44",X"00",X"00",X"F0",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"44",X"00",
		X"00",X"78",X"00",X"81",X"03",X"C0",X"89",X"02",X"B2",X"9A",X"81",X"00",X"78",X"80",X"41",X"00",
		X"03",X"48",X"00",X"80",X"45",X"00",X"03",X"48",X"00",X"80",X"48",X"00",X"02",X"D0",X"00",X"80",
		X"45",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",
		X"00",X"81",X"03",X"C0",X"8A",X"89",X"02",X"B2",X"C9",X"81",X"01",X"E0",X"80",X"34",X"00",X"03",
		X"C0",X"00",X"80",X"3E",X"00",X"03",X"48",X"00",X"80",X"42",X"00",X"00",X"F0",X"00",X"80",X"41",
		X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",
		X"81",X"03",X"C0",X"8A",X"81",X"00",X"F0",X"80",X"4A",X"00",X"03",X"C0",X"00",X"80",X"45",X"00",
		X"01",X"E0",X"00",X"80",X"42",X"00",X"00",X"F0",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",
		X"44",X"00",X"00",X"78",X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"01",X"68",
		X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",
		X"81",X"00",X"F0",X"80",X"4E",X"00",X"03",X"C0",X"00",X"80",X"4A",X"00",X"01",X"E0",X"00",X"80",
		X"48",X"00",X"01",X"68",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"78",
		X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"F0",X"00",X"80",X"4E",X"00",
		X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",X"54",X"00",X"03",
		X"C0",X"00",X"80",X"48",X"00",X"04",X"B0",X"00",X"80",X"46",X"00",X"00",X"F0",X"00",X"80",X"44",
		X"00",X"00",X"F0",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",X"00",
		X"81",X"03",X"C0",X"80",X"44",X"00",X"00",X"F0",X"00",X"80",X"4A",X"00",X"00",X"F0",X"00",X"80",
		X"4D",X"00",X"00",X"F0",X"00",X"80",X"44",X"00",X"00",X"F0",X"00",X"80",X"4A",X"00",X"00",X"F0",
		X"00",X"80",X"44",X"00",X"00",X"F0",X"00",X"80",X"3E",X"00",X"00",X"F0",X"00",X"80",X"4A",X"00",
		X"00",X"F0",X"00",X"80",X"54",X"00",X"01",X"E0",X"00",X"80",X"51",X"00",X"00",X"78",X"00",X"80",
		X"4E",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",
		X"00",X"81",X"03",X"C0",X"89",X"04",X"B3",X"E8",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",
		X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",
		X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",
		X"CF",X"8B",X"0A",X"80",X"44",X"00",X"04",X"38",X"00",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",
		X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",X"00",X"78",
		X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",
		X"9A",X"CF",X"8B",X"0A",X"80",X"44",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"8A",X"89",X"02",
		X"B4",X"52",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"5A",X"00",X"00",X"78",X"00",
		X"80",X"5A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"5A",X"00",X"00",X"78",X"00",X"80",
		X"5A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"4A",X"00",
		X"04",X"38",X"00",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"5A",X"00",X"00",X"78",
		X"00",X"80",X"5A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"5A",X"00",X"00",X"78",X"00",
		X"80",X"5A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"4A",
		X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"8A",X"89",X"02",X"B4",X"BC",X"88",X"9C",X"55",X"8B",
		X"0A",X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"44",X"00",X"04",X"38",X"00",X"88",X"9C",X"55",
		X"8B",X"0A",X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",
		X"00",X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"44",X"00",X"00",X"78",X"00",X"81",X"03",
		X"C0",X"8A",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"5A",X"00",X"00",X"78",X"00",
		X"80",X"5A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"5A",X"00",X"00",X"78",X"00",X"80",
		X"5A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"4A",X"00",
		X"04",X"38",X"00",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"59",X"00",X"00",X"78",
		X"00",X"80",X"59",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"59",X"00",X"00",X"78",X"00",
		X"80",X"59",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"4D",
		X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",
		X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"58",
		X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",
		X"8B",X"0A",X"80",X"4A",X"00",X"04",X"38",X"00",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",
		X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",
		X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",
		X"CF",X"8B",X"0A",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"88",X"9C",X"55",X"8B",
		X"0A",X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"44",X"00",X"04",X"38",X"00",X"88",X"9C",X"55",
		X"8B",X"0A",X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",
		X"00",X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"44",X"00",X"00",X"78",X"00",X"81",X"03",
		X"C0",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",
		X"58",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"58",X"00",X"00",X"78",X"00",X"80",X"58",
		X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"4A",X"00",X"04",
		X"38",X"00",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"55",X"00",X"00",X"78",X"00",
		X"80",X"55",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"55",X"00",X"00",X"78",X"00",X"80",
		X"55",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"4A",X"00",
		X"04",X"38",X"00",X"88",X"9A",X"CF",X"8B",X"03",X"8A",X"88",X"9A",X"CF",X"89",X"00",X"B6",X"C0",
		X"89",X"03",X"B6",X"C4",X"80",X"2A",X"00",X"03",X"C0",X"00",X"80",X"3D",X"00",X"03",X"C0",X"00",
		X"80",X"4A",X"00",X"02",X"D0",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",
		X"78",X"00",X"81",X"03",X"C0",X"8A",X"81",X"01",X"E0",X"80",X"4A",X"00",X"03",X"C0",X"00",X"80",
		X"42",X"00",X"01",X"E0",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",
		X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"F0",X"00",X"80",X"3A",X"00",
		X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"81",
		X"03",X"C0",X"89",X"02",X"B7",X"26",X"80",X"3E",X"00",X"03",X"48",X"00",X"80",X"41",X"00",X"03",
		X"48",X"00",X"80",X"45",X"00",X"01",X"68",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"41",
		X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"F0",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",
		X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"8A",
		X"89",X"02",X"B7",X"64",X"80",X"2A",X"00",X"03",X"C0",X"00",X"80",X"3D",X"00",X"03",X"C0",X"00",
		X"80",X"4A",X"00",X"02",X"D0",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",
		X"78",X"00",X"81",X"03",X"C0",X"8A",X"80",X"48",X"00",X"01",X"E0",X"00",X"80",X"45",X"00",X"01",
		X"E0",X"00",X"80",X"42",X"00",X"01",X"E0",X"00",X"80",X"3E",X"00",X"01",X"E0",X"00",X"80",X"3D",
		X"00",X"01",X"E0",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",
		X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",
		X"4D",X"00",X"01",X"E0",X"00",X"80",X"4A",X"00",X"01",X"E0",X"00",X"80",X"48",X"00",X"01",X"E0",
		X"00",X"80",X"44",X"00",X"01",X"E0",X"00",X"80",X"41",X"00",X"01",X"E0",X"00",X"80",X"49",X"00",
		X"00",X"78",X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",X"45",X"00",X"00",X"78",X"00",X"80",
		X"41",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"81",X"01",X"E0",X"80",X"4A",X"00",X"03",X"C0",
		X"00",X"80",X"42",X"00",X"01",X"E0",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",
		X"00",X"78",X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"F0",X"00",X"80",
		X"3A",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",
		X"00",X"81",X"03",X"C0",X"81",X"00",X"78",X"80",X"3A",X"00",X"00",X"F0",X"00",X"80",X"3D",X"00",
		X"00",X"F0",X"00",X"80",X"3E",X"00",X"00",X"F0",X"00",X"80",X"41",X"00",X"00",X"F0",X"00",X"80",
		X"44",X"00",X"00",X"F0",X"00",X"80",X"3A",X"00",X"00",X"F0",X"00",X"80",X"38",X"00",X"00",X"F0",
		X"00",X"80",X"35",X"00",X"00",X"F0",X"00",X"80",X"3A",X"00",X"00",X"F0",X"00",X"80",X"3E",X"00",
		X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",
		X"3A",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"89",X"04",
		X"B8",X"92",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"4A",X"00",X"00",X"78",X"00",
		X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",
		X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"3A",X"00",
		X"04",X"38",X"00",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"4A",X"00",X"00",X"78",
		X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"4A",X"00",X"00",X"78",X"00",
		X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"3A",
		X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"8A",X"89",X"02",X"B8",X"FC",X"88",X"9C",X"55",X"8B",
		X"0A",X"81",X"00",X"78",X"80",X"51",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"80",X"51",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"41",X"00",X"04",X"38",X"00",X"88",X"9C",X"55",
		X"8B",X"0A",X"81",X"00",X"78",X"80",X"51",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",
		X"00",X"81",X"00",X"78",X"80",X"51",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"41",X"00",X"00",X"78",X"00",X"81",X"03",
		X"C0",X"8A",X"89",X"02",X"B9",X"66",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"4A",
		X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"4A",X"00",
		X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",
		X"0A",X"80",X"3A",X"00",X"04",X"38",X"00",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",
		X"4A",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"4A",
		X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",
		X"8B",X"0A",X"80",X"3A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"8A",X"88",X"9C",X"55",X"8B",
		X"0A",X"81",X"00",X"78",X"80",X"55",X"00",X"00",X"78",X"00",X"80",X"55",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"80",X"55",X"00",X"00",X"78",X"00",X"80",X"55",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"41",X"00",X"04",X"38",X"00",X"88",X"9C",X"55",
		X"8B",X"0A",X"81",X"00",X"78",X"80",X"54",X"00",X"00",X"78",X"00",X"80",X"54",X"00",X"00",X"78",
		X"00",X"81",X"00",X"78",X"80",X"54",X"00",X"00",X"78",X"00",X"80",X"54",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"44",X"00",X"00",X"78",X"00",X"81",X"03",
		X"C0",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"52",X"00",X"00",X"78",X"00",X"80",
		X"52",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"52",X"00",X"00",X"78",X"00",X"80",X"52",
		X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"42",X"00",X"04",
		X"38",X"00",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"51",X"00",X"00",X"78",X"00",
		X"80",X"51",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"51",X"00",X"00",X"78",X"00",X"80",
		X"51",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"41",X"00",
		X"00",X"78",X"00",X"81",X"03",X"C0",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",X"4A",
		X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"4A",X"00",
		X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",X"8B",
		X"0A",X"80",X"3A",X"00",X"04",X"38",X"00",X"88",X"9C",X"55",X"8B",X"0A",X"81",X"00",X"78",X"80",
		X"4A",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"4A",
		X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"88",X"9A",X"CF",
		X"8B",X"0A",X"80",X"3A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"88",X"9C",X"55",X"8B",X"0A",
		X"81",X"00",X"78",X"80",X"54",X"00",X"00",X"78",X"00",X"80",X"54",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"80",X"54",X"00",X"00",X"78",X"00",X"80",X"54",X"00",X"00",X"78",X"00",X"81",X"00",
		X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"54",X"00",X"04",X"38",X"00",X"88",X"9C",X"55",X"8B",
		X"0A",X"81",X"00",X"78",X"80",X"51",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"80",X"51",X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"88",X"9A",X"CF",X"8B",X"0A",X"80",X"54",X"00",X"04",X"38",X"00",X"88",X"9A",X"CF",
		X"8B",X"03",X"8A",X"88",X"9C",X"3B",X"89",X"04",X"BB",X"6A",X"81",X"2D",X"00",X"8A",X"81",X"00",
		X"1E",X"8F",X"AD",X"5F",X"88",X"9B",X"03",X"89",X"00",X"BB",X"7B",X"89",X"04",X"BB",X"7F",X"8C",
		X"00",X"00",X"80",X"1A",X"00",X"01",X"E0",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",
		X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",
		X"8C",X"00",X"00",X"83",X"00",X"F0",X"80",X"1A",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"00",
		X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"1A",
		X"00",X"00",X"78",X"00",X"8C",X"00",X"00",X"83",X"00",X"78",X"80",X"1A",X"00",X"00",X"78",X"00",
		X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",
		X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"26",X"00",X"00",X"78",X"00",X"80",X"1A",
		X"00",X"00",X"78",X"00",X"8C",X"00",X"00",X"81",X"03",X"C0",X"8A",X"89",X"02",X"BB",X"FF",X"8C",
		X"00",X"00",X"80",X"15",X"00",X"00",X"F0",X"00",X"80",X"15",X"00",X"00",X"F0",X"00",X"80",X"21",
		X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"1E",X"00",X"00",X"78",X"00",
		X"80",X"18",X"00",X"00",X"78",X"00",X"8C",X"00",X"00",X"83",X"00",X"F0",X"80",X"18",X"00",X"00",
		X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"80",X"24",
		X"00",X"00",X"78",X"00",X"80",X"1E",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",
		X"8C",X"00",X"00",X"83",X"00",X"78",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"29",X"00",X"00",
		X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"80",X"21",
		X"00",X"00",X"78",X"00",X"80",X"1E",X"00",X"00",X"78",X"00",X"80",X"11",X"00",X"00",X"78",X"00",
		X"8C",X"00",X"00",X"81",X"03",X"C0",X"8A",X"89",X"02",X"BC",X"8B",X"8C",X"00",X"00",X"80",X"1A",
		X"00",X"01",X"E0",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"8C",X"00",X"00",X"83",
		X"00",X"F0",X"80",X"1A",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",
		X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",
		X"8C",X"00",X"00",X"83",X"00",X"78",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",
		X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"28",
		X"00",X"00",X"78",X"00",X"80",X"26",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",
		X"8C",X"00",X"00",X"81",X"03",X"C0",X"8A",X"8C",X"00",X"00",X"80",X"25",X"00",X"00",X"F0",X"00",
		X"80",X"25",X"00",X"00",X"F0",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",
		X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"8C",X"00",
		X"01",X"83",X"00",X"F0",X"80",X"25",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",
		X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",
		X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"8C",X"00",X"00",X"83",X"00",X"F0",X"80",X"24",
		X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",
		X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",
		X"78",X"00",X"8C",X"00",X"00",X"81",X"03",X"C0",X"8C",X"00",X"00",X"80",X"22",X"00",X"00",X"F0",
		X"00",X"80",X"22",X"00",X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",
		X"00",X"78",X"00",X"80",X"26",X"00",X"00",X"78",X"00",X"80",X"22",X"00",X"00",X"78",X"00",X"8C",
		X"00",X"02",X"83",X"00",X"78",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"26",X"00",
		X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"8C",X"00",X"00",X"83",X"00",X"F0",X"80",
		X"21",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"21",X"00",
		X"00",X"78",X"00",X"8C",X"00",X"00",X"81",X"03",X"C0",X"8C",X"00",X"00",X"80",X"1A",X"00",X"01",
		X"E0",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",
		X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"8C",X"00",X"00",X"83",X"00",X"F0",
		X"80",X"1A",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",
		X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"8C",X"00",
		X"00",X"83",X"00",X"78",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",
		X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",
		X"78",X"00",X"80",X"26",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"8C",X"00",
		X"00",X"81",X"03",X"C0",X"8C",X"00",X"00",X"80",X"28",X"00",X"00",X"F0",X"00",X"80",X"28",X"00",
		X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",
		X"2A",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"26",X"00",X"00",X"78",
		X"00",X"8C",X"00",X"00",X"83",X"00",X"F0",X"80",X"26",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",
		X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",
		X"1A",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"8C",X"00",X"01",X"83",X"00",
		X"78",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",
		X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",
		X"2A",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"8C",X"00",X"00",X"83",X"02",
		X"D0",X"80",X"22",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"8A",X"BF",X"2E",
		X"BF",X"39",X"C1",X"AE",X"C4",X"35",X"C6",X"F8",X"C7",X"32",X"9D",X"F5",X"9F",X"79",X"88",X"9B",
		X"1D",X"89",X"00",X"BF",X"35",X"8F",X"A6",X"9A",X"8A",X"88",X"9B",X"37",X"89",X"00",X"BF",X"40",
		X"89",X"02",X"BF",X"44",X"81",X"02",X"58",X"80",X"54",X"00",X"02",X"D0",X"00",X"80",X"48",X"00",
		X"01",X"68",X"00",X"80",X"51",X"00",X"01",X"E0",X"00",X"80",X"4E",X"00",X"01",X"E0",X"00",X"80",
		X"4A",X"00",X"01",X"E0",X"00",X"80",X"51",X"00",X"01",X"68",X"00",X"80",X"44",X"00",X"00",X"F0",
		X"00",X"80",X"4E",X"00",X"01",X"E0",X"00",X"80",X"4A",X"00",X"00",X"F0",X"00",X"80",X"48",X"00",
		X"01",X"68",X"00",X"80",X"4E",X"00",X"00",X"F0",X"00",X"80",X"41",X"00",X"01",X"68",X"00",X"80",
		X"4A",X"00",X"00",X"78",X"00",X"80",X"48",X"00",X"01",X"68",X"00",X"80",X"44",X"00",X"01",X"68",
		X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"38",X"00",
		X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"90",X"88",X"9B",X"51",X"81",X"00",X"F0",
		X"81",X"00",X"78",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"01",X"E0",X"00",X"88",
		X"9B",X"37",X"8A",X"81",X"02",X"58",X"80",X"51",X"00",X"02",X"D0",X"00",X"80",X"4E",X"00",X"01",
		X"68",X"00",X"80",X"4D",X"00",X"01",X"E0",X"00",X"80",X"4E",X"00",X"01",X"E0",X"00",X"80",X"4A",
		X"00",X"01",X"E0",X"00",X"80",X"41",X"00",X"01",X"68",X"00",X"80",X"4E",X"00",X"00",X"F0",X"00",
		X"80",X"48",X"00",X"01",X"E0",X"00",X"80",X"45",X"00",X"00",X"F0",X"00",X"80",X"41",X"00",X"01",
		X"68",X"00",X"80",X"48",X"00",X"00",X"F0",X"00",X"80",X"45",X"00",X"01",X"68",X"00",X"80",X"49",
		X"00",X"00",X"78",X"00",X"80",X"48",X"00",X"01",X"68",X"00",X"80",X"45",X"00",X"01",X"68",X"00",
		X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",
		X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"88",X"9B",X"51",X"81",X"00",X"F0",X"80",X"51",
		X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"F0",X"00",X"80",X"41",X"00",X"00",X"F0",X"00",
		X"80",X"3E",X"00",X"00",X"78",X"00",X"88",X"9B",X"37",X"8F",X"BF",X"44",X"88",X"9B",X"51",X"81",
		X"00",X"F0",X"80",X"4A",X"00",X"00",X"F0",X"00",X"80",X"5A",X"00",X"00",X"78",X"00",X"80",X"54",
		X"00",X"00",X"78",X"00",X"80",X"5D",X"00",X"00",X"F0",X"00",X"88",X"9B",X"37",X"81",X"02",X"58",
		X"80",X"52",X"00",X"02",X"D0",X"00",X"80",X"4E",X"00",X"01",X"68",X"00",X"80",X"45",X"00",X"01",
		X"E0",X"00",X"80",X"42",X"00",X"01",X"E0",X"00",X"80",X"4D",X"00",X"01",X"E0",X"00",X"80",X"51",
		X"00",X"01",X"68",X"00",X"80",X"4E",X"00",X"00",X"F0",X"00",X"80",X"4D",X"00",X"01",X"E0",X"00",
		X"80",X"4E",X"00",X"00",X"F0",X"00",X"80",X"49",X"00",X"01",X"68",X"00",X"80",X"4A",X"00",X"00",
		X"F0",X"00",X"80",X"42",X"00",X"01",X"68",X"00",X"80",X"4D",X"00",X"00",X"78",X"00",X"80",X"4E",
		X"00",X"01",X"68",X"00",X"80",X"52",X"00",X"01",X"68",X"00",X"80",X"51",X"00",X"00",X"78",X"00",
		X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",
		X"78",X"00",X"88",X"9B",X"51",X"81",X"00",X"F0",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"48",
		X"00",X"00",X"78",X"00",X"80",X"4A",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"01",X"68",X"00",
		X"88",X"9B",X"37",X"81",X"02",X"58",X"80",X"54",X"00",X"02",X"D0",X"00",X"80",X"48",X"00",X"01",
		X"68",X"00",X"80",X"51",X"00",X"01",X"E0",X"00",X"80",X"4E",X"00",X"01",X"E0",X"00",X"80",X"4A",
		X"00",X"01",X"E0",X"00",X"80",X"51",X"00",X"01",X"68",X"00",X"80",X"44",X"00",X"00",X"F0",X"00",
		X"80",X"4E",X"00",X"01",X"E0",X"00",X"80",X"4A",X"00",X"00",X"F0",X"00",X"80",X"48",X"00",X"01",
		X"68",X"00",X"80",X"46",X"00",X"00",X"F0",X"00",X"80",X"4A",X"00",X"01",X"68",X"00",X"80",X"45",
		X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"01",X"68",X"00",X"80",X"3E",X"00",X"01",X"68",X"00",
		X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",
		X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"88",X"9B",X"51",X"81",X"00",X"F0",X"80",X"54",
		X"00",X"00",X"78",X"00",X"80",X"51",X"00",X"02",X"58",X"00",X"88",X"9B",X"37",X"8A",X"88",X"9B",
		X"37",X"89",X"00",X"C1",X"B5",X"89",X"02",X"C1",X"B9",X"81",X"01",X"E0",X"80",X"44",X"00",X"01",
		X"E0",X"00",X"80",X"3E",X"00",X"01",X"E0",X"00",X"80",X"41",X"00",X"02",X"58",X"00",X"80",X"38",
		X"00",X"01",X"E0",X"00",X"80",X"41",X"00",X"01",X"E0",X"00",X"80",X"3A",X"00",X"01",X"68",X"00",
		X"80",X"3E",X"00",X"01",X"E0",X"00",X"80",X"36",X"00",X"01",X"E0",X"00",X"80",X"3E",X"00",X"00",
		X"F0",X"00",X"80",X"38",X"00",X"01",X"68",X"00",X"80",X"3A",X"00",X"00",X"F0",X"00",X"80",X"31",
		X"00",X"00",X"F0",X"00",X"80",X"3A",X"00",X"00",X"F0",X"00",X"80",X"34",X"00",X"00",X"F0",X"00",
		X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"38",X"00",X"00",
		X"78",X"00",X"80",X"36",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"34",
		X"00",X"00",X"78",X"00",X"90",X"88",X"9B",X"51",X"81",X"00",X"F0",X"81",X"00",X"50",X"80",X"38",
		X"00",X"00",X"50",X"00",X"80",X"3A",X"00",X"00",X"50",X"00",X"80",X"3D",X"00",X"01",X"E0",X"00",
		X"88",X"9B",X"37",X"8A",X"81",X"01",X"E0",X"80",X"3A",X"00",X"01",X"E0",X"00",X"80",X"38",X"00",
		X"01",X"E0",X"00",X"80",X"34",X"00",X"02",X"58",X"00",X"80",X"3A",X"00",X"01",X"E0",X"00",X"80",
		X"38",X"00",X"01",X"E0",X"00",X"80",X"35",X"00",X"01",X"68",X"00",X"80",X"34",X"00",X"01",X"E0",
		X"00",X"80",X"35",X"00",X"01",X"E0",X"00",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"2E",X"00",
		X"01",X"68",X"00",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"00",X"F0",X"00",X"80",
		X"34",X"00",X"00",X"F0",X"00",X"80",X"35",X"00",X"00",X"F0",X"00",X"80",X"38",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"38",X"00",
		X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"88",
		X"9B",X"51",X"81",X"00",X"F0",X"81",X"00",X"50",X"80",X"4E",X"00",X"00",X"F0",X"00",X"80",X"41",
		X"00",X"00",X"50",X"00",X"80",X"48",X"00",X"01",X"40",X"00",X"88",X"9B",X"37",X"8F",X"C1",X"B9",
		X"88",X"9B",X"51",X"81",X"00",X"F0",X"81",X"00",X"50",X"80",X"48",X"00",X"00",X"50",X"00",X"80",
		X"4A",X"00",X"02",X"30",X"00",X"88",X"9B",X"37",X"81",X"01",X"E0",X"80",X"3E",X"00",X"01",X"E0",
		X"00",X"80",X"42",X"00",X"01",X"E0",X"00",X"80",X"41",X"00",X"02",X"58",X"00",X"80",X"3E",X"00",
		X"01",X"E0",X"00",X"80",X"3D",X"00",X"01",X"E0",X"00",X"80",X"3A",X"00",X"01",X"68",X"00",X"80",
		X"38",X"00",X"01",X"E0",X"00",X"80",X"34",X"00",X"01",X"E0",X"00",X"80",X"32",X"00",X"00",X"F0",
		X"00",X"80",X"3A",X"00",X"01",X"68",X"00",X"80",X"3E",X"00",X"00",X"F0",X"00",X"80",X"36",X"00",
		X"00",X"F0",X"00",X"80",X"34",X"00",X"00",X"F0",X"00",X"80",X"32",X"00",X"00",X"F0",X"00",X"80",
		X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"31",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",
		X"00",X"78",X"00",X"88",X"9B",X"51",X"81",X"00",X"F0",X"81",X"00",X"50",X"80",X"2E",X"00",X"00",
		X"50",X"00",X"80",X"31",X"00",X"01",X"E0",X"00",X"80",X"3A",X"00",X"00",X"50",X"00",X"88",X"9B",
		X"37",X"81",X"01",X"E0",X"80",X"44",X"00",X"01",X"E0",X"00",X"80",X"3E",X"00",X"01",X"E0",X"00",
		X"80",X"41",X"00",X"02",X"58",X"00",X"80",X"38",X"00",X"01",X"E0",X"00",X"80",X"41",X"00",X"01",
		X"E0",X"00",X"80",X"3A",X"00",X"01",X"68",X"00",X"80",X"3E",X"00",X"01",X"E0",X"00",X"80",X"34",
		X"00",X"01",X"E0",X"00",X"80",X"32",X"00",X"00",X"F0",X"00",X"80",X"31",X"00",X"01",X"68",X"00",
		X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"00",
		X"F0",X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2D",
		X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",
		X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"88",X"9B",X"51",X"81",
		X"00",X"F0",X"81",X"01",X"40",X"80",X"54",X"00",X"00",X"50",X"00",X"80",X"51",X"00",X"01",X"40",
		X"00",X"88",X"9B",X"37",X"8A",X"88",X"9B",X"37",X"89",X"00",X"C4",X"3C",X"89",X"02",X"C4",X"40",
		X"80",X"2A",X"00",X"02",X"58",X"00",X"80",X"2E",X"00",X"01",X"E0",X"00",X"80",X"31",X"00",X"01",
		X"68",X"00",X"80",X"2E",X"00",X"01",X"E0",X"00",X"80",X"31",X"00",X"01",X"E0",X"00",X"80",X"32",
		X"00",X"01",X"E0",X"00",X"80",X"34",X"00",X"01",X"68",X"00",X"80",X"38",X"00",X"01",X"68",X"00",
		X"80",X"3A",X"00",X"01",X"68",X"00",X"80",X"38",X"00",X"01",X"68",X"00",X"80",X"3A",X"00",X"01",
		X"68",X"00",X"80",X"34",X"00",X"00",X"F0",X"00",X"80",X"32",X"00",X"00",X"F0",X"00",X"80",X"31",
		X"00",X"01",X"68",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"F0",X"00",
		X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2D",
		X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"90",X"88",X"9B",X"51",X"81",X"01",
		X"2C",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"02",X"1C",X"00",X"88",X"9B",X"37",
		X"8A",X"80",X"21",X"00",X"02",X"58",X"00",X"80",X"25",X"00",X"01",X"E0",X"00",X"80",X"28",X"00",
		X"01",X"68",X"00",X"80",X"25",X"00",X"01",X"E0",X"00",X"80",X"28",X"00",X"01",X"E0",X"00",X"80",
		X"29",X"00",X"01",X"E0",X"00",X"80",X"2A",X"00",X"01",X"68",X"00",X"80",X"2E",X"00",X"01",X"68",
		X"00",X"80",X"31",X"00",X"01",X"68",X"00",X"80",X"2E",X"00",X"01",X"68",X"00",X"80",X"31",X"00",
		X"01",X"68",X"00",X"80",X"2A",X"00",X"00",X"F0",X"00",X"80",X"29",X"00",X"00",X"F0",X"00",X"80",
		X"28",X"00",X"01",X"68",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"F0",
		X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",
		X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"80",
		X"24",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"51",X"81",X"02",
		X"94",X"80",X"44",X"00",X"00",X"3C",X"00",X"80",X"41",X"00",X"00",X"F0",X"00",X"88",X"9B",X"37",
		X"8F",X"C4",X"40",X"88",X"9B",X"51",X"81",X"00",X"F0",X"80",X"44",X"00",X"00",X"78",X"00",X"80",
		X"38",X"00",X"02",X"1C",X"00",X"80",X"44",X"00",X"00",X"3C",X"00",X"88",X"9B",X"37",X"80",X"25",
		X"00",X"02",X"58",X"00",X"80",X"2E",X"00",X"01",X"E0",X"00",X"80",X"32",X"00",X"01",X"68",X"00",
		X"80",X"2E",X"00",X"01",X"E0",X"00",X"80",X"2D",X"00",X"01",X"E0",X"00",X"80",X"28",X"00",X"01",
		X"E0",X"00",X"80",X"24",X"00",X"01",X"68",X"00",X"80",X"2A",X"00",X"01",X"68",X"00",X"80",X"28",
		X"00",X"01",X"68",X"00",X"80",X"2E",X"00",X"01",X"68",X"00",X"80",X"2A",X"00",X"01",X"68",X"00",
		X"80",X"22",X"00",X"00",X"F0",X"00",X"80",X"32",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"01",
		X"68",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"26",X"00",X"00",X"F0",X"00",X"80",X"2E",
		X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",
		X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"88",X"9B",X"51",X"81",X"00",X"F0",X"81",X"00",
		X"3C",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"31",X"00",
		X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",
		X"28",X"00",X"00",X"3C",X"00",X"88",X"9B",X"37",X"80",X"2A",X"00",X"02",X"58",X"00",X"80",X"2E",
		X"00",X"01",X"E0",X"00",X"80",X"31",X"00",X"01",X"68",X"00",X"80",X"2E",X"00",X"01",X"E0",X"00",
		X"80",X"31",X"00",X"01",X"E0",X"00",X"80",X"32",X"00",X"01",X"E0",X"00",X"80",X"34",X"00",X"01",
		X"68",X"00",X"80",X"38",X"00",X"01",X"68",X"00",X"80",X"3A",X"00",X"01",X"68",X"00",X"80",X"3A",
		X"00",X"01",X"68",X"00",X"80",X"2A",X"00",X"01",X"68",X"00",X"80",X"3A",X"00",X"00",X"F0",X"00",
		X"80",X"2A",X"00",X"00",X"F0",X"00",X"80",X"3A",X"00",X"01",X"68",X"00",X"80",X"2A",X"00",X"00",
		X"78",X"00",X"80",X"3A",X"00",X"00",X"F0",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"3A",
		X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",
		X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",
		X"78",X"00",X"88",X"9B",X"51",X"81",X"03",X"0C",X"80",X"42",X"00",X"00",X"78",X"00",X"80",X"41",
		X"00",X"00",X"3C",X"00",X"88",X"9B",X"37",X"8A",X"89",X"00",X"C6",X"FC",X"89",X"21",X"C7",X"00",
		X"8C",X"01",X"00",X"81",X"03",X"C0",X"8A",X"8C",X"01",X"01",X"81",X"03",X"C0",X"89",X"03",X"C7",
		X"11",X"8C",X"01",X"00",X"81",X"03",X"C0",X"8A",X"8C",X"01",X"02",X"81",X"03",X"C0",X"89",X"0A",
		X"C7",X"22",X"8C",X"01",X"00",X"81",X"03",X"C0",X"8A",X"8A",X"89",X"00",X"C7",X"2E",X"81",X"25",
		X"80",X"8A",X"88",X"9B",X"03",X"89",X"00",X"C7",X"39",X"89",X"02",X"C7",X"3D",X"80",X"1A",X"00",
		X"03",X"48",X"00",X"80",X"24",X"00",X"03",X"C0",X"00",X"80",X"28",X"00",X"03",X"C0",X"00",X"80",
		X"31",X"00",X"03",X"C0",X"00",X"80",X"34",X"00",X"02",X"58",X"00",X"80",X"32",X"00",X"01",X"E0",
		X"00",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",
		X"00",X"F0",X"00",X"80",X"28",X"00",X"00",X"F0",X"00",X"80",X"1A",X"00",X"01",X"E0",X"00",X"80",
		X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",
		X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"90",X"8A",X"80",X"21",X"00",X"03",
		X"48",X"00",X"80",X"2E",X"00",X"01",X"E0",X"00",X"80",X"31",X"00",X"01",X"68",X"00",X"80",X"35",
		X"00",X"00",X"F0",X"00",X"80",X"29",X"00",X"02",X"D0",X"00",X"80",X"21",X"00",X"00",X"78",X"00",
		X"80",X"28",X"00",X"01",X"E0",X"00",X"80",X"31",X"00",X"01",X"68",X"00",X"80",X"35",X"00",X"00",
		X"F0",X"00",X"80",X"25",X"00",X"00",X"F0",X"00",X"80",X"21",X"00",X"01",X"E0",X"00",X"80",X"2E",
		X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"01",X"E0",X"00",X"80",X"35",X"00",X"01",X"68",X"00",
		X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",
		X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",
		X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",
		X"80",X"21",X"00",X"01",X"68",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",
		X"F0",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",
		X"00",X"00",X"78",X"00",X"8F",X"C7",X"3D",X"80",X"25",X"00",X"03",X"48",X"00",X"80",X"32",X"00",
		X"01",X"E0",X"00",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",
		X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"01",X"68",
		X"00",X"80",X"2D",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",
		X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",
		X"31",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",
		X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",
		X"00",X"78",X"00",X"80",X"22",X"00",X"03",X"C0",X"00",X"80",X"2E",X"00",X"01",X"E0",X"00",X"80",
		X"2D",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"26",X"00",X"00",X"78",
		X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"22",X"00",X"00",X"78",X"00",X"80",X"21",X"00",
		X"00",X"F0",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"F0",X"00",X"80",
		X"26",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"F0",
		X"00",X"80",X"32",X"00",X"00",X"F0",X"00",X"80",X"3A",X"00",X"00",X"F0",X"00",X"80",X"3E",X"00",
		X"00",X"F0",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"03",X"48",X"00",X"80",
		X"34",X"00",X"03",X"C0",X"00",X"80",X"3D",X"00",X"03",X"C0",X"00",X"80",X"3A",X"00",X"01",X"E0",
		X"00",X"80",X"38",X"00",X"00",X"F0",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"38",X"00",
		X"00",X"78",X"00",X"80",X"39",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"01",X"68",X"00",X"80",
		X"1E",X"00",X"01",X"E0",X"00",X"80",X"21",X"00",X"01",X"E0",X"00",X"80",X"22",X"00",X"01",X"E0",
		X"00",X"80",X"24",X"00",X"00",X"F0",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"1E",X"00",
		X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"F0",X"00",X"80",X"1E",X"00",X"00",X"78",X"00",X"80",
		X"1A",X"00",X"00",X"78",X"00",X"80",X"14",X"00",X"01",X"68",X"00",X"81",X"02",X"D0",X"8A",X"A6",
		X"93",X"C9",X"9F",X"C9",X"D9",X"C9",X"EB",X"C9",X"FD",X"CE",X"A1",X"9D",X"F5",X"9F",X"79",X"89",
		X"00",X"C9",X"A3",X"89",X"21",X"C9",X"A7",X"8C",X"02",X"00",X"81",X"03",X"C0",X"8A",X"8C",X"02",
		X"01",X"81",X"03",X"C0",X"89",X"03",X"C9",X"B8",X"8C",X"02",X"00",X"81",X"03",X"C0",X"8A",X"8C",
		X"02",X"02",X"81",X"03",X"C0",X"89",X"0A",X"C9",X"C9",X"8C",X"02",X"00",X"81",X"03",X"C0",X"8A",
		X"8A",X"89",X"00",X"C9",X"D5",X"81",X"1E",X"00",X"8A",X"88",X"9D",X"8D",X"94",X"16",X"04",X"94",
		X"17",X"04",X"94",X"18",X"04",X"94",X"19",X"04",X"8F",X"CA",X"00",X"88",X"9D",X"8D",X"94",X"16",
		X"03",X"94",X"17",X"03",X"94",X"18",X"03",X"94",X"19",X"03",X"8F",X"CA",X"00",X"88",X"9D",X"8D",
		X"89",X"00",X"CA",X"04",X"80",X"1A",X"00",X"01",X"E0",X"00",X"80",X"1A",X"00",X"01",X"68",X"00",
		X"80",X"18",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",
		X"1E",X"00",X"01",X"E0",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"1D",
		X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"18",X"00",X"00",X"78",X"00",X"81",X"00",X"78",
		X"80",X"18",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",
		X"1A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",X"24",X"00",X"01",X"E0",X"00",X"80",X"24",
		X"00",X"01",X"68",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"80",X"28",X"00",X"01",X"E0",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"80",X"26",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"21",X"00",X"00",X"78",
		X"00",X"81",X"00",X"78",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",
		X"81",X"00",X"78",X"80",X"1A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",X"1A",X"00",X"00",
		X"F0",X"00",X"80",X"1D",X"00",X"00",X"F0",X"00",X"80",X"1E",X"00",X"00",X"F0",X"00",X"80",X"1D",
		X"00",X"01",X"68",X"00",X"80",X"1E",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"F0",X"00",
		X"80",X"1E",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"18",X"00",X"00",X"F0",X"00",X"80",
		X"1A",X"00",X"00",X"F0",X"00",X"80",X"1D",X"00",X"00",X"F0",X"00",X"80",X"1E",X"00",X"00",X"F0",
		X"00",X"80",X"21",X"00",X"01",X"68",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"25",X"00",
		X"00",X"F0",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"2A",X"00",X"00",
		X"F0",X"00",X"80",X"24",X"00",X"00",X"F0",X"00",X"80",X"26",X"00",X"00",X"F0",X"00",X"80",X"28",
		X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"01",X"68",X"00",X"80",X"28",X"00",X"00",X"78",X"00",
		X"80",X"26",X"00",X"00",X"F0",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"26",X"00",X"00",
		X"78",X"00",X"80",X"21",X"00",X"00",X"F0",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"81",X"00",
		X"78",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"1D",X"00",X"00",X"78",X"00",
		X"80",X"1E",X"00",X"00",X"F0",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",
		X"21",X"00",X"01",X"E0",X"00",X"80",X"21",X"00",X"01",X"68",X"00",X"80",X"1E",X"00",X"00",X"78",
		X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"25",X"00",X"01",X"E0",X"00",
		X"80",X"28",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"24",X"00",X"00",X"78",X"00",X"81",
		X"00",X"78",X"80",X"1E",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"1E",X"00",X"00",X"78",
		X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"21",X"00",X"00",X"78",X"00",
		X"81",X"03",X"C0",X"80",X"21",X"00",X"00",X"F0",X"00",X"89",X"03",X"CB",X"CD",X"80",X"31",X"00",
		X"00",X"78",X"00",X"8A",X"81",X"00",X"78",X"80",X"21",X"00",X"01",X"E0",X"00",X"80",X"31",X"00",
		X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",
		X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"F0",X"00",X"80",X"21",X"00",X"00",X"78",
		X"00",X"81",X"00",X"78",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"00",X"F0",X"00",
		X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",
		X"1A",X"00",X"01",X"E0",X"00",X"80",X"1A",X"00",X"01",X"68",X"00",X"80",X"18",X"00",X"00",X"78",
		X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"1D",X"00",
		X"01",X"68",X"00",X"80",X"1E",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",
		X"1D",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"F0",X"00",X"80",X"1E",X"00",X"00",X"78",
		X"00",X"80",X"1D",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"1E",X"00",
		X"00",X"78",X"00",X"80",X"1D",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"81",
		X"03",X"C0",X"80",X"1A",X"00",X"00",X"F0",X"00",X"80",X"18",X"00",X"00",X"78",X"00",X"80",X"1A",
		X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"1D",X"00",X"00",X"78",X"00",
		X"80",X"1E",X"00",X"01",X"68",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"1D",X"00",X"00",
		X"78",X"00",X"80",X"18",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"1E",
		X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"1D",X"00",X"00",X"78",X"00",
		X"80",X"1E",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",
		X"78",X"00",X"80",X"1D",X"00",X"00",X"F0",X"00",X"80",X"1E",X"00",X"00",X"78",X"00",X"80",X"1D",
		X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",X"2A",X"00",
		X"00",X"F0",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",
		X"2E",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"2E",X"00",X"01",X"E0",X"00",X"80",X"31",
		X"00",X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",
		X"80",X"2A",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"00",X"F0",X"00",X"80",X"28",X"00",X"00",
		X"F0",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"1D",X"00",X"00",X"78",X"00",X"80",X"24",
		X"00",X"00",X"F0",X"00",X"81",X"03",X"C0",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",
		X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"F0",X"00",X"80",
		X"2E",X"00",X"01",X"E0",X"00",X"80",X"2D",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",X"00",X"F0",
		X"00",X"80",X"26",X"00",X"00",X"78",X"00",X"80",X"29",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",
		X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"00",X"F0",X"00",X"80",
		X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",X"2A",
		X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",
		X"80",X"34",X"00",X"01",X"68",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"28",
		X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",
		X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"24",
		X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"80",X"34",X"00",
		X"00",X"F0",X"00",X"89",X"03",X"CE",X"27",X"80",X"34",X"00",X"00",X"78",X"00",X"8A",X"81",X"00",
		X"78",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",
		X"00",X"78",X"00",X"80",X"36",X"00",X"01",X"68",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",
		X"2E",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",
		X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",
		X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",
		X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"80",X"24",
		X"00",X"01",X"E0",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"8A",X"88",X"9B",X"03",X"89",X"00",X"CE",X"A8",X"89",X"04",X"CE",X"AC",X"89",X"05",X"CE",X"B0",
		X"80",X"1A",X"00",X"00",X"B4",X"00",X"81",X"01",X"2C",X"8A",X"80",X"2A",X"00",X"00",X"F0",X"00",
		X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"90",
		X"8A",X"89",X"02",X"CE",X"D5",X"89",X"05",X"CE",X"D9",X"80",X"21",X"00",X"00",X"B4",X"00",X"81",
		X"01",X"2C",X"8A",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",
		X"21",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"8A",X"89",X"02",X"CE",X"FD",X"8F",X"CE",X"AC",
		X"8A",X"89",X"04",X"CF",X"05",X"80",X"25",X"00",X"00",X"B4",X"00",X"81",X"01",X"2C",X"8A",X"80",
		X"24",X"00",X"00",X"B4",X"00",X"81",X"01",X"2C",X"80",X"34",X"00",X"00",X"F0",X"00",X"80",X"24",
		X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"89",X"04",X"CF",
		X"31",X"80",X"22",X"00",X"00",X"B4",X"00",X"81",X"01",X"2C",X"8A",X"80",X"21",X"00",X"00",X"B4",
		X"00",X"81",X"01",X"2C",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"21",X"00",X"00",X"78",X"00",
		X"80",X"21",X"00",X"00",X"78",X"00",X"81",X"03",X"C0",X"8F",X"CE",X"AC",X"89",X"02",X"CF",X"60",
		X"80",X"28",X"00",X"00",X"B4",X"00",X"81",X"01",X"2C",X"8A",X"89",X"02",X"CF",X"6E",X"80",X"26",
		X"00",X"00",X"B4",X"00",X"81",X"01",X"2C",X"8A",X"80",X"25",X"00",X"00",X"B4",X"00",X"81",X"01",
		X"2C",X"80",X"3E",X"00",X"00",X"F0",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"80",X"24",X"00",
		X"00",X"78",X"00",X"81",X"03",X"C0",X"8A",X"D4",X"F2",X"D5",X"24",X"D5",X"32",X"D5",X"CC",X"D6",
		X"A1",X"D7",X"8E",X"9D",X"F5",X"9F",X"79",X"80",X"1A",X"00",X"00",X"78",X"00",X"89",X"04",X"CF",
		X"B1",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"8A",X"80",X"2A",
		X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"18",X"00",X"00",X"78",X"00",
		X"80",X"1A",X"00",X"01",X"E0",X"00",X"90",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"24",X"00",
		X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",
		X"2D",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",
		X"00",X"80",X"1E",X"00",X"00",X"78",X"00",X"90",X"89",X"02",X"D0",X"0C",X"80",X"28",X"00",X"00",
		X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"24",
		X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",
		X"8A",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"24",X"00",
		X"00",X"78",X"00",X"80",X"1E",X"00",X"00",X"78",X"00",X"90",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",
		X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",
		X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",
		X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"36",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"38",
		X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"90",X"80",X"2D",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"90",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2D",
		X"00",X"00",X"78",X"00",X"90",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",
		X"00",X"90",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"90",X"80",
		X"34",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"90",X"80",X"38",X"00",X"00",
		X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"90",X"80",X"38",X"00",X"00",X"78",X"00",X"80",
		X"3A",X"00",X"00",X"78",X"00",X"90",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",
		X"78",X"00",X"90",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",
		X"31",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"90",X"80",X"2A",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"3E",
		X"00",X"00",X"78",X"00",X"80",X"4D",X"00",X"00",X"78",X"00",X"80",X"4E",X"00",X"00",X"78",X"00",
		X"80",X"46",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"90",X"80",X"4E",X"00",
		X"00",X"78",X"00",X"80",X"48",X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",
		X"4A",X"00",X"00",X"78",X"00",X"90",X"89",X"02",X"D1",X"7A",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",
		X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"8A",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",
		X"3A",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"90",X"80",X"21",
		X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",
		X"80",X"28",X"00",X"00",X"78",X"00",X"90",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",
		X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"90",
		X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"31",
		X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",
		X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",
		X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"31",
		X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",
		X"90",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"31",X"00",
		X"00",X"78",X"00",X"90",X"80",X"3E",X"00",X"00",X"78",X"00",X"89",X"02",X"D2",X"6E",X"80",X"41",
		X"00",X"00",X"78",X"00",X"8A",X"90",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",
		X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"90",X"80",X"45",X"00",X"00",X"78",X"00",X"80",
		X"3E",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"90",X"80",X"35",X"00",X"00",
		X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"32",
		X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"90",X"80",X"25",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",
		X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",
		X"3D",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3C",X"00",X"00",X"78",
		X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",
		X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"80",
		X"35",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"78",X"00",X"90",X"80",X"3E",X"00",X"00",
		X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"90",X"80",X"32",X"00",X"00",X"78",X"00",X"80",
		X"35",X"00",X"00",X"78",X"00",X"90",X"80",X"24",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"2D",
		X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",
		X"80",X"24",X"00",X"00",X"78",X"00",X"90",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",
		X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"90",
		X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",
		X"78",X"00",X"80",X"26",X"00",X"00",X"78",X"00",X"80",X"24",X"00",X"00",X"78",X"00",X"90",X"80",
		X"34",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"36",X"00",X"00",X"78",
		X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",
		X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"90",
		X"80",X"54",X"00",X"00",X"78",X"00",X"80",X"4D",X"00",X"00",X"78",X"00",X"80",X"46",X"00",X"00",
		X"78",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",
		X"00",X"00",X"78",X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",
		X"90",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"90",X"80",X"3D",
		X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"90",X"80",X"3E",X"00",X"00",X"78",
		X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"42",X"00",
		X"00",X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"90",
		X"80",X"46",X"00",X"00",X"78",X"00",X"80",X"42",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",
		X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"3A",
		X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",X"36",X"00",X"00",X"78",X"00",
		X"90",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"39",X"00",
		X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"90",X"80",X"32",X"00",X"00",X"78",X"00",
		X"80",X"31",X"00",X"00",X"78",X"00",X"90",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"32",X"00",
		X"00",X"78",X"00",X"90",X"80",X"36",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",
		X"90",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"36",X"00",X"00",X"78",X"00",X"90",X"80",X"3E",
		X"00",X"00",X"78",X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"90",X"80",X"3D",X"00",X"00",X"78",
		X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"90",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"39",
		X"00",X"00",X"78",X"00",X"90",X"80",X"39",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",
		X"00",X"90",X"89",X"00",X"D4",X"F6",X"89",X"21",X"D4",X"FA",X"8C",X"03",X"00",X"81",X"03",X"C0",
		X"8A",X"8C",X"03",X"01",X"81",X"03",X"C0",X"89",X"03",X"D5",X"0B",X"8C",X"03",X"00",X"81",X"03",
		X"C0",X"8A",X"8C",X"03",X"02",X"81",X"03",X"C0",X"89",X"0A",X"D5",X"1C",X"8C",X"03",X"00",X"81",
		X"03",X"C0",X"8A",X"8A",X"88",X"9D",X"A7",X"94",X"19",X"01",X"89",X"00",X"D5",X"2E",X"8F",X"A6",
		X"9A",X"8A",X"89",X"00",X"D5",X"36",X"88",X"9D",X"DB",X"89",X"02",X"D5",X"3D",X"94",X"21",X"1F",
		X"97",X"21",X"FF",X"00",X"7B",X"1F",X"89",X"02",X"D5",X"4A",X"8F",X"D0",X"4A",X"8A",X"8F",X"D1",
		X"2C",X"8F",X"D1",X"76",X"81",X"03",X"C0",X"8A",X"94",X"19",X"04",X"89",X"03",X"D5",X"5F",X"8F",
		X"D1",X"F0",X"96",X"19",X"01",X"8A",X"94",X"19",X"02",X"8F",X"D1",X"D7",X"81",X"00",X"78",X"8F",
		X"D2",X"51",X"81",X"03",X"C0",X"94",X"21",X"1F",X"97",X"21",X"FF",X"00",X"7B",X"1F",X"89",X"02",
		X"D5",X"82",X"8F",X"D0",X"4A",X"8A",X"8F",X"D1",X"2C",X"8F",X"D1",X"76",X"81",X"03",X"C0",X"8F",
		X"D2",X"BB",X"8F",X"D3",X"36",X"8F",X"D3",X"67",X"81",X"01",X"E0",X"8F",X"D4",X"40",X"8F",X"D4",
		X"40",X"94",X"19",X"04",X"8F",X"D1",X"BE",X"94",X"19",X"02",X"81",X"00",X"78",X"8F",X"D2",X"51",
		X"81",X"03",X"C0",X"94",X"19",X"04",X"81",X"01",X"E0",X"8F",X"CF",X"A7",X"8F",X"CF",X"A7",X"94",
		X"19",X"02",X"8F",X"CF",X"A7",X"8F",X"D1",X"13",X"81",X"03",X"C0",X"8A",X"89",X"00",X"D5",X"D0",
		X"88",X"9D",X"DB",X"89",X"02",X"D5",X"D7",X"94",X"21",X"18",X"89",X"08",X"D5",X"DE",X"8F",X"D0",
		X"AB",X"8F",X"D0",X"AB",X"96",X"21",X"03",X"8A",X"8F",X"D0",X"4A",X"8F",X"D0",X"C5",X"8F",X"D0",
		X"EC",X"8F",X"D0",X"C5",X"8F",X"D0",X"F9",X"81",X"03",X"C0",X"8A",X"89",X"02",X"D5",X"FF",X"94",
		X"19",X"01",X"89",X"02",X"D6",X"06",X"81",X"00",X"78",X"8F",X"D2",X"76",X"8A",X"94",X"19",X"02",
		X"8F",X"D2",X"51",X"81",X"00",X"78",X"8F",X"D1",X"BE",X"8A",X"8F",X"D1",X"F0",X"8F",X"D1",X"BE",
		X"8F",X"D1",X"D7",X"81",X"03",X"C0",X"94",X"21",X"18",X"89",X"08",X"D6",X"2D",X"8F",X"D0",X"AB",
		X"8F",X"D0",X"AB",X"96",X"21",X"03",X"8A",X"8F",X"D0",X"4A",X"8F",X"D0",X"C5",X"8F",X"D0",X"EC",
		X"8F",X"D0",X"C5",X"8F",X"D0",X"F9",X"81",X"03",X"C0",X"81",X"00",X"78",X"89",X"03",X"D6",X"50",
		X"8F",X"D2",X"9C",X"8A",X"89",X"02",X"D6",X"58",X"8F",X"D3",X"80",X"8A",X"8F",X"D3",X"67",X"8F",
		X"D4",X"01",X"94",X"19",X"01",X"8F",X"D4",X"40",X"8F",X"D4",X"71",X"8F",X"D4",X"71",X"94",X"19",
		X"02",X"8F",X"D2",X"51",X"81",X"00",X"F0",X"8F",X"D2",X"64",X"81",X"03",X"C0",X"89",X"02",X"D6",
		X"81",X"8F",X"CF",X"D7",X"8A",X"8F",X"D0",X"08",X"94",X"19",X"04",X"8F",X"CF",X"A7",X"94",X"19",
		X"02",X"8F",X"D0",X"AB",X"8F",X"D0",X"C5",X"8F",X"D0",X"F9",X"8F",X"D0",X"EC",X"81",X"03",X"C0",
		X"8A",X"88",X"9D",X"DB",X"89",X"00",X"D6",X"A8",X"89",X"02",X"D6",X"AC",X"89",X"02",X"D6",X"B0",
		X"8F",X"CF",X"A7",X"8A",X"81",X"00",X"78",X"89",X"08",X"D6",X"BB",X"8F",X"D0",X"B8",X"8A",X"8F",
		X"D0",X"EC",X"81",X"00",X"78",X"89",X"02",X"D6",X"C9",X"8F",X"D0",X"F9",X"8A",X"81",X"03",X"C0",
		X"8A",X"81",X"00",X"F0",X"89",X"03",X"D6",X"D8",X"8F",X"D1",X"BE",X"81",X"00",X"78",X"8A",X"8F",
		X"D2",X"51",X"81",X"00",X"78",X"8F",X"D2",X"76",X"89",X"02",X"D6",X"EC",X"81",X"00",X"78",X"8F",
		X"D2",X"64",X"8A",X"94",X"19",X"04",X"89",X"02",X"D6",X"FA",X"8F",X"D1",X"BE",X"8A",X"94",X"19",
		X"02",X"8F",X"D1",X"F0",X"81",X"03",X"C0",X"89",X"02",X"D7",X"0B",X"8F",X"CF",X"A7",X"8A",X"81",
		X"00",X"78",X"89",X"08",X"D7",X"16",X"8F",X"D0",X"B8",X"8A",X"8F",X"D0",X"EC",X"81",X"00",X"78",
		X"89",X"02",X"D7",X"24",X"8F",X"D0",X"F9",X"8A",X"81",X"03",X"C0",X"81",X"00",X"78",X"94",X"19",
		X"01",X"89",X"03",X"D7",X"35",X"8F",X"D3",X"1C",X"8F",X"D3",X"29",X"8A",X"8F",X"D2",X"89",X"94",
		X"19",X"02",X"89",X"02",X"D7",X"46",X"8F",X"D3",X"36",X"8A",X"94",X"19",X"00",X"89",X"03",X"D7",
		X"51",X"8F",X"D4",X"1B",X"95",X"19",X"01",X"8A",X"89",X"02",X"D7",X"5C",X"94",X"19",X"02",X"8F",
		X"D2",X"76",X"8A",X"81",X"03",X"C0",X"89",X"02",X"D7",X"6A",X"8F",X"D0",X"08",X"8A",X"94",X"19",
		X"00",X"89",X"08",X"D7",X"75",X"8F",X"D0",X"F9",X"95",X"19",X"01",X"8A",X"89",X"04",X"D7",X"80",
		X"8F",X"D0",X"EC",X"96",X"19",X"02",X"8A",X"81",X"03",X"C0",X"94",X"19",X"02",X"8A",X"88",X"9B",
		X"03",X"89",X"00",X"D7",X"95",X"89",X"02",X"D7",X"99",X"80",X"1A",X"00",X"02",X"58",X"00",X"80",
		X"24",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"01",X"E0",
		X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",X"24",X"00",
		X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"26",X"00",X"01",X"E0",X"00",X"80",
		X"2E",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",
		X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"F0",X"00",X"89",X"02",X"D7",
		X"F1",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"8A",X"80",X"2A",
		X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",
		X"90",X"80",X"24",X"00",X"01",X"68",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"22",X"00",
		X"00",X"F0",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"01",X"E0",X"00",X"80",
		X"2A",X"00",X"00",X"78",X"00",X"80",X"20",X"00",X"00",X"F0",X"00",X"80",X"1A",X"00",X"00",X"78",
		X"00",X"80",X"1E",X"00",X"00",X"F0",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",
		X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"80",
		X"22",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"F0",
		X"00",X"81",X"03",X"48",X"90",X"8A",X"80",X"21",X"00",X"02",X"58",X"00",X"80",X"2A",X"00",X"00",
		X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"01",X"E0",X"00",X"80",X"31",
		X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",
		X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"F0",X"00",X"80",X"31",X"00",X"00",
		X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"F0",X"00",X"80",X"31",
		X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"2C",X"00",X"01",X"68",X"00",
		X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",
		X"78",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"2A",
		X"00",X"00",X"F0",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",
		X"80",X"29",X"00",X"00",X"F0",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",
		X"78",X"00",X"80",X"28",X"00",X"00",X"F0",X"00",X"80",X"35",X"00",X"00",X"78",X"00",X"80",X"34",
		X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",
		X"80",X"29",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",
		X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"F0",X"00",X"80",X"28",
		X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",
		X"80",X"21",X"00",X"00",X"F0",X"00",X"81",X"03",X"48",X"8F",X"D7",X"99",X"8F",X"D8",X"11",X"80",
		X"25",X"00",X"02",X"58",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"35",X"00",X"00",X"78",
		X"00",X"80",X"38",X"00",X"01",X"E0",X"00",X"80",X"35",X"00",X"00",X"F0",X"00",X"80",X"34",X"00",
		X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",
		X"24",X"00",X"02",X"58",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",
		X"00",X"80",X"38",X"00",X"00",X"F0",X"00",X"80",X"36",X"00",X"00",X"F0",X"00",X"80",X"34",X"00",
		X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",
		X"22",X"00",X"02",X"D0",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"00",X"F0",X"00",X"80",X"2A",X"00",
		X"00",X"F0",X"00",X"80",X"1E",X"00",X"00",X"F0",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",
		X"21",X"00",X"00",X"78",X"00",X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",
		X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",
		X"00",X"78",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"F0",X"00",X"81",
		X"03",X"48",X"8F",X"D7",X"99",X"80",X"24",X"00",X"01",X"68",X"00",X"80",X"2A",X"00",X"00",X"78",
		X"00",X"80",X"2E",X"00",X"00",X"F0",X"00",X"80",X"1A",X"00",X"00",X"78",X"00",X"80",X"28",X"00",
		X"01",X"E0",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"26",X"00",X"00",X"F0",X"00",X"80",
		X"1A",X"00",X"00",X"78",X"00",X"80",X"25",X"00",X"00",X"F0",X"00",X"80",X"21",X"00",X"00",X"78",
		X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",
		X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"22",X"00",X"00",X"78",X"00",X"80",
		X"24",X"00",X"00",X"F0",X"00",X"81",X"03",X"48",X"8A",X"80",X"44",X"00",X"00",X"78",X"00",X"80",
		X"34",X"00",X"00",X"78",X"00",X"80",X"3D",X"00",X"00",X"78",X"00",X"80",X"44",X"00",X"00",X"78",
		X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"38",X"00",
		X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"90",X"88",X"9B",X"03",X"80",X"24",X"00",
		X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"32",X"00",X"00",X"78",X"00",X"80",
		X"31",X"00",X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",
		X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"90",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"3A",
		X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",
		X"80",X"31",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"38",X"00",X"00",
		X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"90",X"88",X"9B",X"03",X"80",X"21",X"00",X"00",
		X"78",X"00",X"80",X"22",X"00",X"00",X"78",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"24",
		X"00",X"00",X"F0",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"80",X"21",X"00",X"00",X"78",X"00",
		X"80",X"1E",X"00",X"00",X"78",X"00",X"90",X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"3C",X"00",
		X"80",X"21",X"00",X"00",X"3C",X"00",X"81",X"01",X"E0",X"88",X"9B",X"D3",X"80",X"28",X"00",X"00",
		X"78",X"00",X"80",X"28",X"00",X"00",X"78",X"00",X"88",X"9B",X"85",X"80",X"21",X"00",X"00",X"3C",
		X"00",X"80",X"21",X"00",X"00",X"3C",X"00",X"90",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",
		X"FF",X"00",X"07",X"08",X"80",X"21",X"00",X"00",X"3C",X"00",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"07",X"08",X"80",X"21",X"00",X"00",X"3C",X"00",X"88",X"9A",X"9B",X"94",X"12",X"21",X"97",
		X"12",X"FF",X"00",X"0F",X"10",X"80",X"21",X"00",X"00",X"F0",X"00",X"94",X"12",X"21",X"97",X"12",
		X"FF",X"00",X"0F",X"10",X"80",X"21",X"00",X"00",X"F0",X"00",X"88",X"9B",X"B9",X"94",X"12",X"30",
		X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",X"03",X"80",X"30",X"00",X"00",
		X"78",X"00",X"94",X"12",X"30",X"97",X"12",X"FF",X"00",X"07",X"08",X"97",X"12",X"FF",X"00",X"28",
		X"03",X"80",X"30",X"00",X"00",X"78",X"00",X"88",X"9B",X"6B",X"94",X"12",X"21",X"97",X"12",X"FF",
		X"00",X"07",X"08",X"80",X"21",X"00",X"00",X"3C",X"00",X"94",X"12",X"21",X"97",X"12",X"FF",X"00",
		X"07",X"08",X"80",X"21",X"00",X"00",X"3C",X"00",X"90",X"89",X"00",X"DC",X"1D",X"81",X"1E",X"00",
		X"8A",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"31",X"DC",X"39",X"DC",X"3F",X"DC",
		X"45",X"88",X"9A",X"B5",X"8F",X"DA",X"99",X"8E",X"01",X"8F",X"DA",X"CA",X"8F",X"DC",X"19",X"8F",
		X"DB",X"57",X"8F",X"DC",X"19",X"8F",X"DB",X"88",X"8F",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",
		X"19",X"DC",X"19",X"DC",X"5B",X"DC",X"39",X"DC",X"3F",X"DC",X"45",X"88",X"9B",X"1D",X"8F",X"DA",
		X"99",X"8E",X"02",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"73",X"DC",X"39",X"DC",
		X"3F",X"DC",X"45",X"88",X"9A",X"B5",X"8F",X"DA",X"99",X"8E",X"03",X"DC",X"19",X"DC",X"19",X"DC",
		X"19",X"DC",X"19",X"DC",X"8B",X"DC",X"39",X"DC",X"3F",X"DC",X"45",X"88",X"9D",X"A7",X"94",X"19",
		X"01",X"8F",X"DA",X"99",X"8E",X"04",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"A6",
		X"DC",X"AE",X"DC",X"3F",X"DC",X"45",X"88",X"9A",X"B5",X"8F",X"DA",X"F8",X"8E",X"01",X"8F",X"DB",
		X"29",X"8F",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"C4",X"DC",X"AE",
		X"DC",X"3F",X"DC",X"45",X"88",X"9B",X"1D",X"8F",X"DA",X"F8",X"8E",X"02",X"DC",X"19",X"DC",X"19",
		X"DC",X"19",X"DC",X"19",X"DC",X"DC",X"DC",X"AE",X"DC",X"3F",X"DC",X"45",X"88",X"9A",X"B5",X"8F",
		X"DA",X"F8",X"8E",X"03",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"19",X"DC",X"F4",X"DC",X"AE",
		X"DC",X"3F",X"DC",X"45",X"88",X"9D",X"A7",X"8F",X"DA",X"F8",X"8E",X"04",X"0F",X"DD",X"05",X"DD",
		X"0B",X"DD",X"11",X"DD",X"17",X"81",X"03",X"FC",X"8F",X"DD",X"17",X"81",X"02",X"94",X"8F",X"DD",
		X"17",X"81",X"01",X"A4",X"8F",X"DD",X"17",X"88",X"9A",X"CF",X"80",X"2A",X"00",X"00",X"3C",X"00",
		X"80",X"31",X"00",X"00",X"3C",X"00",X"80",X"34",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"00",
		X"3C",X"00",X"80",X"36",X"00",X"00",X"3C",X"00",X"80",X"34",X"00",X"00",X"3C",X"00",X"80",X"44",
		X"00",X"01",X"68",X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",X"80",X"46",X"00",X"00",X"3C",X"00",
		X"80",X"44",X"00",X"00",X"3C",X"00",X"80",X"50",X"00",X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",
		X"3C",X"00",X"80",X"44",X"00",X"00",X"3C",X"00",X"80",X"3A",X"00",X"02",X"D0",X"00",X"92",X"0F",
		X"DD",X"78",X"DD",X"97",X"DD",X"B6",X"DD",X"D5",X"88",X"9C",X"21",X"80",X"3A",X"00",X"00",X"B4",
		X"00",X"81",X"00",X"3C",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",
		X"80",X"44",X"00",X"03",X"C0",X"00",X"92",X"88",X"9C",X"07",X"80",X"34",X"00",X"00",X"B4",X"00",
		X"81",X"00",X"3C",X"80",X"34",X"00",X"00",X"78",X"00",X"80",X"34",X"00",X"00",X"78",X"00",X"80",
		X"3A",X"00",X"03",X"C0",X"00",X"92",X"88",X"9C",X"07",X"80",X"2A",X"00",X"00",X"B4",X"00",X"81",
		X"00",X"3C",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"00",X"78",X"00",X"80",X"2D",
		X"00",X"03",X"C0",X"00",X"92",X"88",X"9B",X"03",X"80",X"2A",X"00",X"00",X"B4",X"00",X"81",X"00",
		X"3C",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"3A",X"00",X"00",X"78",X"00",X"80",X"2A",X"00",
		X"03",X"C0",X"00",X"92",X"0F",X"DD",X"FD",X"DD",X"FD",X"DD",X"FD",X"DD",X"FD",X"88",X"9A",X"CF",
		X"94",X"12",X"44",X"97",X"12",X"01",X"00",X"25",X"10",X"80",X"44",X"00",X"02",X"58",X"00",X"88",
		X"9B",X"51",X"94",X"2D",X"0A",X"80",X"44",X"00",X"03",X"C0",X"00",X"92",X"0F",X"DE",X"25",X"DE",
		X"4E",X"DE",X"5B",X"DE",X"68",X"88",X"9A",X"CF",X"89",X"04",X"DE",X"2C",X"94",X"12",X"24",X"97",
		X"12",X"01",X"00",X"06",X"30",X"80",X"24",X"00",X"01",X"2C",X"00",X"8B",X"08",X"8A",X"88",X"9B",
		X"51",X"94",X"2D",X"09",X"8B",X"08",X"90",X"80",X"34",X"00",X"03",X"C0",X"00",X"92",X"81",X"00",
		X"3C",X"8F",X"DE",X"25",X"80",X"2D",X"00",X"03",X"C0",X"00",X"92",X"81",X"00",X"8C",X"8F",X"DE",
		X"25",X"80",X"2A",X"00",X"03",X"C0",X"00",X"92",X"81",X"00",X"E1",X"8F",X"DE",X"25",X"80",X"1A",
		X"00",X"03",X"C0",X"00",X"92",X"0F",X"DE",X"7E",X"DE",X"D0",X"DE",X"D6",X"DE",X"DC",X"88",X"9A",
		X"CF",X"80",X"2A",X"00",X"00",X"5A",X"00",X"80",X"31",X"00",X"00",X"5A",X"00",X"80",X"34",X"00",
		X"00",X"5A",X"00",X"80",X"38",X"00",X"00",X"5A",X"00",X"80",X"34",X"00",X"00",X"5A",X"00",X"80",
		X"3A",X"00",X"00",X"5A",X"00",X"80",X"38",X"00",X"00",X"5A",X"00",X"80",X"41",X"00",X"00",X"5A",
		X"00",X"80",X"3E",X"00",X"00",X"5A",X"00",X"80",X"3A",X"00",X"00",X"5A",X"00",X"80",X"38",X"00",
		X"00",X"5A",X"00",X"80",X"41",X"00",X"00",X"2D",X"00",X"80",X"44",X"00",X"02",X"58",X"00",X"92",
		X"81",X"00",X"3C",X"8F",X"DE",X"7E",X"81",X"00",X"C8",X"8F",X"DE",X"7E",X"81",X"01",X"08",X"8F",
		X"DE",X"7E",X"07",X"DE",X"E9",X"DE",X"E9",X"DE",X"E9",X"88",X"9C",X"BD",X"94",X"12",X"34",X"97",
		X"12",X"FF",X"00",X"18",X"0A",X"80",X"34",X"00",X"00",X"F0",X"00",X"92",X"07",X"DF",X"03",X"DF",
		X"03",X"DF",X"03",X"88",X"9C",X"F1",X"94",X"12",X"34",X"97",X"12",X"FF",X"00",X"78",X"03",X"80",
		X"34",X"00",X"01",X"68",X"00",X"92",X"07",X"DF",X"1D",X"DF",X"1D",X"DF",X"1D",X"88",X"9D",X"0B",
		X"80",X"34",X"00",X"01",X"68",X"00",X"92",X"3F",X"DF",X"34",X"DF",X"41",X"DF",X"4E",X"DF",X"5B",
		X"DF",X"34",X"DF",X"34",X"88",X"9A",X"67",X"94",X"35",X"0A",X"80",X"04",X"00",X"05",X"A0",X"00",
		X"92",X"88",X"9A",X"67",X"94",X"35",X"0B",X"80",X"15",X"00",X"04",X"B0",X"00",X"92",X"88",X"9A",
		X"67",X"94",X"35",X"0C",X"80",X"26",X"00",X"03",X"FC",X"00",X"92",X"88",X"9A",X"67",X"94",X"35",
		X"0D",X"80",X"38",X"00",X"03",X"84",X"00",X"92",X"FF",X"DF",X"AD",X"DF",X"BA",X"DF",X"C7",X"DF",
		X"D4",X"DF",X"AD",X"DF",X"BA",X"DF",X"C7",X"DF",X"D4",X"88",X"9A",X"67",X"94",X"35",X"0E",X"80",
		X"24",X"00",X"01",X"A4",X"00",X"92",X"88",X"9A",X"67",X"94",X"35",X"0E",X"80",X"22",X"00",X"01",
		X"E0",X"00",X"92",X"88",X"9A",X"67",X"94",X"35",X"0D",X"80",X"15",X"00",X"02",X"58",X"00",X"92",
		X"88",X"9A",X"67",X"94",X"35",X"0C",X"80",X"12",X"00",X"03",X"48",X"00",X"92",X"88",X"9A",X"67",
		X"94",X"35",X"0B",X"80",X"2D",X"00",X"04",X"74",X"00",X"92",X"88",X"9A",X"67",X"94",X"35",X"0A",
		X"80",X"1E",X"00",X"05",X"DC",X"00",X"92",X"88",X"9A",X"67",X"94",X"35",X"09",X"80",X"15",X"00",
		X"07",X"80",X"00",X"92",X"88",X"9A",X"67",X"94",X"35",X"09",X"80",X"04",X"00",X"09",X"60",X"00",
		X"92",X"FF",X"E0",X"C2",X"E0",X"A9",X"E0",X"99",X"E0",X"89",X"E0",X"69",X"E0",X"41",X"E0",X"1D",
		X"DF",X"F2",X"88",X"9A",X"67",X"80",X"2D",X"00",X"00",X"F0",X"00",X"80",X"2D",X"00",X"01",X"E0",
		X"00",X"80",X"2D",X"00",X"01",X"E0",X"00",X"80",X"2D",X"00",X"00",X"78",X"00",X"80",X"2D",X"00",
		X"00",X"78",X"00",X"94",X"35",X"0E",X"80",X"2D",X"00",X"01",X"E0",X"00",X"92",X"88",X"9A",X"67",
		X"81",X"00",X"5A",X"80",X"2C",X"00",X"02",X"58",X"00",X"94",X"35",X"11",X"89",X"07",X"E0",X"30",
		X"80",X"1C",X"00",X"00",X"3C",X"00",X"8A",X"94",X"35",X"0D",X"80",X"1C",X"00",X"02",X"D0",X"00",
		X"92",X"88",X"9A",X"67",X"81",X"00",X"96",X"80",X"14",X"00",X"04",X"B0",X"00",X"80",X"14",X"00",
		X"00",X"B4",X"00",X"80",X"14",X"00",X"00",X"78",X"00",X"80",X"14",X"00",X"00",X"78",X"00",X"94",
		X"35",X"0A",X"80",X"14",X"00",X"04",X"B0",X"00",X"92",X"88",X"9A",X"CF",X"89",X"08",X"E0",X"70",
		X"94",X"12",X"14",X"80",X"14",X"00",X"00",X"0F",X"00",X"89",X"0F",X"E0",X"7D",X"95",X"12",X"03",
		X"83",X"00",X"0F",X"8A",X"8B",X"04",X"8A",X"90",X"92",X"88",X"9A",X"67",X"81",X"00",X"78",X"80",
		X"04",X"00",X"00",X"F0",X"00",X"8F",X"E0",X"69",X"92",X"88",X"9A",X"67",X"81",X"00",X"B4",X"80",
		X"04",X"00",X"00",X"F0",X"00",X"8F",X"E0",X"69",X"92",X"81",X"00",X"3C",X"8F",X"E0",X"69",X"88",
		X"9A",X"67",X"80",X"05",X"00",X"00",X"F0",X"00",X"94",X"35",X"07",X"80",X"05",X"00",X"09",X"60",
		X"00",X"92",X"81",X"00",X"96",X"8F",X"E0",X"69",X"88",X"9A",X"67",X"80",X"04",X"00",X"00",X"F0",
		X"00",X"94",X"35",X"07",X"80",X"04",X"00",X"09",X"60",X"00",X"92",X"0F",X"E0",X"E4",X"E0",X"E4",
		X"E0",X"E4",X"E0",X"E4",X"88",X"9C",X"6F",X"80",X"25",X"00",X"00",X"F0",X"00",X"92",X"0F",X"E0",
		X"F7",X"E0",X"F7",X"E0",X"F7",X"E0",X"F7",X"88",X"9C",X"6F",X"80",X"15",X"00",X"02",X"58",X"00",
		X"92",X"0F",X"E1",X"0A",X"E1",X"0A",X"E1",X"0A",X"E1",X"0A",X"88",X"9C",X"A3",X"94",X"12",X"34",
		X"97",X"12",X"01",X"00",X"0B",X"20",X"80",X"34",X"00",X"01",X"68",X"00",X"92",X"0F",X"E1",X"26",
		X"E1",X"26",X"E1",X"42",X"E1",X"68",X"88",X"9C",X"6F",X"94",X"17",X"06",X"97",X"17",X"FF",X"00",
		X"30",X"05",X"94",X"21",X"1F",X"97",X"21",X"FF",X"00",X"07",X"1F",X"80",X"18",X"00",X"00",X"F0",
		X"00",X"92",X"88",X"9B",X"85",X"94",X"1F",X"12",X"94",X"21",X"14",X"94",X"2B",X"0A",X"94",X"2C",
		X"00",X"94",X"2D",X"0D",X"94",X"35",X"0A",X"90",X"94",X"12",X"5E",X"97",X"12",X"FF",X"00",X"07",
		X"20",X"80",X"5E",X"00",X"00",X"F0",X"00",X"92",X"8F",X"E1",X"42",X"94",X"12",X"58",X"97",X"12",
		X"FF",X"00",X"07",X"20",X"80",X"58",X"00",X"00",X"F0",X"00",X"92",X"07",X"E1",X"82",X"E1",X"AE",
		X"E1",X"B4",X"88",X"9B",X"51",X"94",X"41",X"00",X"89",X"05",X"E1",X"8C",X"80",X"44",X"00",X"00",
		X"5A",X"00",X"80",X"2D",X"00",X"00",X"5A",X"00",X"80",X"51",X"00",X"00",X"5A",X"00",X"80",X"3A",
		X"00",X"00",X"5A",X"00",X"80",X"18",X"00",X"00",X"5A",X"00",X"8B",X"07",X"8A",X"92",X"81",X"00",
		X"50",X"8F",X"E1",X"82",X"81",X"00",X"84",X"8F",X"E1",X"82",X"0F",X"E1",X"C3",X"E1",X"C3",X"E1",
		X"C3",X"E1",X"C3",X"88",X"9B",X"9F",X"80",X"44",X"00",X"00",X"B4",X"00",X"92",X"FF",X"E1",X"DE",
		X"E1",X"DE",X"E1",X"DE",X"E1",X"DE",X"E1",X"DE",X"E1",X"DE",X"E1",X"DE",X"E1",X"DE",X"88",X"9A",
		X"81",X"80",X"22",X"00",X"01",X"68",X"00",X"92",X"FF",X"E1",X"F9",X"E1",X"F9",X"E1",X"F9",X"E1",
		X"F9",X"E1",X"F9",X"E1",X"F9",X"E1",X"F9",X"E1",X"F9",X"88",X"9C",X"D7",X"94",X"12",X"2A",X"97",
		X"12",X"01",X"00",X"18",X"0A",X"80",X"2A",X"00",X"00",X"F0",X"00",X"88",X"9C",X"BD",X"94",X"12",
		X"34",X"97",X"12",X"FF",X"00",X"18",X"0A",X"80",X"34",X"00",X"00",X"F0",X"00",X"92",X"0F",X"E2",
		X"27",X"E2",X"27",X"E2",X"27",X"E2",X"27",X"88",X"9D",X"25",X"94",X"13",X"00",X"97",X"13",X"08",
		X"00",X"03",X"1F",X"80",X"54",X"00",X"01",X"2C",X"00",X"92",X"03",X"E2",X"3F",X"E2",X"3F",X"88",
		X"9D",X"3F",X"94",X"1E",X"0C",X"80",X"2A",X"00",X"00",X"F0",X"00",X"92",X"03",X"E2",X"51",X"E2",
		X"7F",X"88",X"9D",X"0B",X"94",X"25",X"0E",X"94",X"19",X"07",X"94",X"35",X"1F",X"80",X"54",X"00",
		X"00",X"F0",X"00",X"81",X"00",X"5A",X"94",X"25",X"1F",X"80",X"4C",X"00",X"00",X"3C",X"00",X"81",
		X"00",X"3C",X"94",X"25",X"0E",X"94",X"35",X"1F",X"80",X"54",X"00",X"01",X"68",X"00",X"92",X"88",
		X"9D",X"0B",X"94",X"25",X"0E",X"94",X"19",X"06",X"94",X"39",X"40",X"94",X"35",X"1F",X"81",X"01",
		X"86",X"80",X"42",X"00",X"01",X"2C",X"00",X"92",X"01",X"E2",X"9B",X"88",X"9B",X"51",X"89",X"02",
		X"E2",X"A2",X"80",X"54",X"00",X"00",X"5A",X"00",X"8A",X"88",X"9B",X"37",X"80",X"54",X"00",X"00",
		X"3C",X"00",X"80",X"3A",X"00",X"00",X"B4",X"00",X"88",X"9D",X"3F",X"8B",X"0A",X"94",X"1E",X"0D",
		X"80",X"44",X"00",X"00",X"F0",X"00",X"92",X"0F",X"E2",X"D0",X"E2",X"FE",X"E3",X"09",X"E3",X"14",
		X"88",X"9D",X"3F",X"94",X"1E",X"0D",X"80",X"2A",X"00",X"00",X"78",X"00",X"88",X"9A",X"CF",X"80",
		X"34",X"00",X"00",X"5A",X"00",X"80",X"3A",X"00",X"00",X"5A",X"00",X"80",X"3D",X"00",X"00",X"5A",
		X"00",X"80",X"44",X"00",X"00",X"5A",X"00",X"80",X"54",X"00",X"01",X"E0",X"00",X"92",X"81",X"00",
		X"B4",X"88",X"9A",X"CF",X"8B",X"06",X"8F",X"E2",X"DF",X"81",X"01",X"2C",X"88",X"9A",X"CF",X"8B",
		X"0C",X"8F",X"E2",X"DF",X"81",X"01",X"7C",X"88",X"9A",X"CF",X"8B",X"12",X"8F",X"E2",X"DF",X"0F",
		X"E3",X"2B",X"E3",X"4A",X"E3",X"55",X"E3",X"60",X"88",X"9B",X"9F",X"80",X"34",X"00",X"00",X"3C",
		X"00",X"80",X"3C",X"00",X"00",X"78",X"00",X"81",X"00",X"F0",X"80",X"3C",X"00",X"00",X"3C",X"00",
		X"80",X"32",X"00",X"00",X"78",X"00",X"81",X"00",X"78",X"92",X"81",X"00",X"0F",X"88",X"9B",X"9F",
		X"8B",X"04",X"8F",X"E3",X"2B",X"81",X"00",X"18",X"88",X"9B",X"9F",X"8B",X"07",X"8F",X"E3",X"2B",
		X"81",X"00",X"28",X"88",X"9B",X"9F",X"8B",X"0B",X"8F",X"E3",X"2B",X"0F",X"E3",X"B6",X"E3",X"A0",
		X"E3",X"8A",X"E3",X"74",X"88",X"9A",X"67",X"81",X"00",X"F0",X"80",X"08",X"00",X"00",X"F0",X"00",
		X"94",X"35",X"08",X"80",X"08",X"00",X"07",X"80",X"00",X"92",X"88",X"9A",X"67",X"81",X"00",X"B4",
		X"80",X"06",X"00",X"00",X"F0",X"00",X"94",X"35",X"08",X"80",X"06",X"00",X"07",X"80",X"00",X"92",
		X"81",X"00",X"3C",X"88",X"9A",X"67",X"80",X"05",X"00",X"00",X"F0",X"00",X"94",X"35",X"07",X"80",
		X"05",X"00",X"0B",X"40",X"00",X"92",X"88",X"9A",X"67",X"80",X"04",X"00",X"00",X"F0",X"00",X"94",
		X"35",X"07",X"80",X"04",X"00",X"0B",X"40",X"00",X"92",X"03",X"E3",X"CE",X"E3",X"FB",X"88",X"9A",
		X"81",X"94",X"20",X"22",X"94",X"21",X"1A",X"80",X"24",X"00",X"00",X"3C",X"00",X"89",X"00",X"E3",
		X"E1",X"94",X"21",X"1A",X"97",X"21",X"FF",X"00",X"03",X"1A",X"83",X"00",X"5A",X"94",X"21",X"00",
		X"97",X"21",X"01",X"00",X"03",X"1A",X"83",X"00",X"5A",X"8A",X"92",X"88",X"9A",X"81",X"94",X"19",
		X"02",X"81",X"00",X"2D",X"8F",X"E3",X"D1",X"0F",X"E4",X"10",X"E4",X"43",X"E4",X"76",X"E4",X"A9",
		X"88",X"9A",X"CF",X"80",X"64",X"00",X"00",X"B4",X"00",X"94",X"12",X"64",X"97",X"12",X"FF",X"00",
		X"08",X"30",X"83",X"02",X"1C",X"88",X"9D",X"59",X"8B",X"05",X"94",X"12",X"2C",X"97",X"12",X"FF",
		X"00",X"0F",X"08",X"97",X"12",X"FF",X"00",X"50",X"03",X"80",X"2C",X"00",X"00",X"F0",X"00",X"83",
		X"01",X"68",X"92",X"88",X"9A",X"CF",X"80",X"4A",X"00",X"00",X"B4",X"00",X"94",X"12",X"4A",X"97",
		X"12",X"FF",X"00",X"13",X"16",X"83",X"02",X"3A",X"88",X"9D",X"59",X"8B",X"09",X"94",X"12",X"2C",
		X"97",X"12",X"FF",X"00",X"0F",X"08",X"97",X"12",X"FF",X"00",X"50",X"03",X"80",X"2C",X"00",X"00",
		X"F0",X"00",X"83",X"01",X"68",X"92",X"88",X"9A",X"CF",X"80",X"18",X"00",X"00",X"B4",X"00",X"94",
		X"12",X"18",X"97",X"12",X"01",X"00",X"0F",X"1C",X"83",X"02",X"44",X"88",X"9D",X"59",X"8B",X"0D",
		X"94",X"12",X"2C",X"97",X"12",X"FF",X"00",X"0F",X"08",X"97",X"12",X"FF",X"00",X"50",X"03",X"80",
		X"2C",X"00",X"00",X"F0",X"00",X"83",X"01",X"68",X"92",X"88",X"9A",X"CF",X"80",X"00",X"00",X"00",
		X"B4",X"00",X"94",X"12",X"00",X"97",X"12",X"01",X"00",X"08",X"34",X"83",X"02",X"49",X"88",X"9D",
		X"59",X"8B",X"10",X"94",X"12",X"2C",X"97",X"12",X"FF",X"00",X"0F",X"08",X"97",X"12",X"FF",X"00",
		X"50",X"03",X"80",X"2C",X"00",X"00",X"F0",X"00",X"83",X"01",X"68",X"92",X"0F",X"E4",X"E5",X"E5",
		X"2B",X"E5",X"36",X"E5",X"41",X"88",X"9A",X"CF",X"80",X"4E",X"00",X"00",X"78",X"00",X"80",X"4A",
		X"00",X"00",X"78",X"00",X"80",X"48",X"00",X"00",X"3C",X"00",X"80",X"4A",X"00",X"00",X"3C",X"00",
		X"80",X"48",X"00",X"00",X"3C",X"00",X"80",X"44",X"00",X"00",X"78",X"00",X"80",X"42",X"00",X"00",
		X"78",X"00",X"80",X"41",X"00",X"00",X"78",X"00",X"80",X"3E",X"00",X"00",X"78",X"00",X"80",X"3A",
		X"00",X"00",X"78",X"00",X"80",X"2A",X"00",X"02",X"D0",X"00",X"92",X"81",X"00",X"96",X"88",X"9A",
		X"CF",X"8B",X"04",X"8F",X"E4",X"E8",X"81",X"00",X"C3",X"88",X"9A",X"CF",X"8B",X"07",X"8F",X"E4",
		X"E8",X"81",X"01",X"14",X"88",X"9A",X"CF",X"8B",X"0A",X"8F",X"E4",X"E8",X"F0",X"E5",X"55",X"E5",
		X"74",X"E5",X"93",X"E5",X"AF",X"88",X"9B",X"51",X"81",X"00",X"D2",X"80",X"5A",X"00",X"00",X"3C",
		X"00",X"80",X"64",X"00",X"01",X"0E",X"00",X"80",X"62",X"00",X"00",X"78",X"00",X"80",X"56",X"00",
		X"01",X"2C",X"00",X"92",X"88",X"9B",X"51",X"80",X"44",X"00",X"00",X"B4",X"00",X"81",X"00",X"B4",
		X"80",X"55",X"00",X"00",X"78",X"00",X"80",X"59",X"00",X"00",X"3C",X"00",X"80",X"31",X"00",X"00",
		X"B4",X"00",X"92",X"88",X"9B",X"ED",X"89",X"04",X"E5",X"9A",X"94",X"12",X"24",X"97",X"12",X"01",
		X"00",X"03",X"20",X"80",X"24",X"00",X"00",X"78",X"00",X"8B",X"04",X"8A",X"8B",X"F0",X"92",X"88",
		X"9B",X"ED",X"8B",X"10",X"89",X"04",X"E5",X"B8",X"94",X"12",X"55",X"97",X"12",X"FF",X"00",X"02",
		X"20",X"80",X"55",X"00",X"00",X"5A",X"00",X"8B",X"FC",X"8A",X"92",X"3F",X"E5",X"D8",X"E5",X"EA",
		X"E5",X"D8",X"E5",X"EA",X"E5",X"D8",X"E5",X"EA",X"88",X"9D",X"3F",X"8B",X"08",X"94",X"22",X"09",
		X"94",X"1E",X"06",X"80",X"24",X"00",X"02",X"58",X"00",X"92",X"88",X"9D",X"3F",X"8B",X"0C",X"81",
		X"00",X"3C",X"8F",X"E5",X"DD",X"01",X"E5",X"F8",X"88",X"9D",X"59",X"94",X"12",X"2C",X"97",X"12",
		X"FF",X"00",X"0F",X"08",X"97",X"12",X"FF",X"00",X"50",X"03",X"80",X"2C",X"00",X"00",X"F0",X"00",
		X"92",X"FF",X"E6",X"22",X"E6",X"3E",X"E6",X"49",X"E6",X"54",X"E6",X"22",X"E6",X"3E",X"E6",X"49",
		X"E6",X"54",X"88",X"9B",X"9F",X"80",X"24",X"00",X"00",X"3C",X"00",X"80",X"2C",X"00",X"00",X"3C",
		X"00",X"80",X"26",X"00",X"00",X"3C",X"00",X"80",X"2E",X"00",X"00",X"78",X"00",X"92",X"88",X"9B",
		X"9F",X"8B",X"02",X"81",X"00",X"12",X"8F",X"E6",X"25",X"88",X"9B",X"9F",X"8B",X"03",X"81",X"00",
		X"14",X"8F",X"E6",X"25",X"88",X"9B",X"9F",X"8B",X"03",X"81",X"00",X"16",X"8F",X"E6",X"25",X"0F",
		X"E6",X"68",X"E6",X"75",X"E6",X"68",X"E6",X"75",X"88",X"9A",X"67",X"94",X"35",X"0E",X"80",X"04",
		X"00",X"02",X"58",X"00",X"92",X"88",X"9A",X"67",X"94",X"35",X"0F",X"80",X"05",X"00",X"01",X"E0",
		X"00",X"92",X"0F",X"E6",X"8B",X"E6",X"B0",X"E6",X"D5",X"E6",X"FA",X"88",X"9A",X"81",X"94",X"12",
		X"41",X"97",X"12",X"FF",X"00",X"0F",X"30",X"97",X"20",X"FF",X"00",X"0B",X"15",X"80",X"41",X"00",
		X"02",X"D0",X"00",X"88",X"9A",X"67",X"94",X"35",X"0E",X"80",X"01",X"00",X"02",X"58",X"00",X"92",
		X"88",X"9A",X"81",X"94",X"12",X"42",X"97",X"12",X"FF",X"00",X"0F",X"30",X"97",X"20",X"FF",X"00",
		X"0B",X"15",X"80",X"42",X"00",X"02",X"D0",X"00",X"88",X"9A",X"67",X"94",X"35",X"0E",X"80",X"02",
		X"00",X"02",X"58",X"00",X"92",X"88",X"9A",X"81",X"94",X"12",X"44",X"97",X"12",X"FF",X"00",X"0F",
		X"30",X"97",X"20",X"FF",X"00",X"0B",X"15",X"80",X"44",X"00",X"02",X"D0",X"00",X"88",X"9A",X"67",
		X"94",X"35",X"0E",X"80",X"04",X"00",X"02",X"58",X"00",X"92",X"88",X"9A",X"81",X"94",X"12",X"45",
		X"97",X"12",X"FF",X"00",X"0F",X"30",X"97",X"20",X"FF",X"00",X"0B",X"15",X"80",X"45",X"00",X"02",
		X"D0",X"00",X"88",X"9A",X"67",X"94",X"35",X"0E",X"80",X"05",X"00",X"02",X"58",X"00",X"92",X"10",
		X"CE",X"07",X"FC",X"CC",X"8A",X"12",X"FD",X"07",X"FD",X"7E",X"80",X"01",X"E7",X"1F",X"80",X"45",
		X"82",X"1F",X"80",X"45",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"10",X"CE",X"07",X"FF",X"8E",X"E7",X"2C",X"48",X"6E",X"96",
		X"80",X"45",X"FF",X"F0",X"FF",X"F0",X"80",X"01",X"82",X"1F",X"FF",X"F0",X"82",X"1F",X"80",X"45");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
