library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity joust2_bg_sound_bank_b is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of joust2_bg_sound_bank_b is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"DD",X"19",X"0A",X"17",X"26",X"0A",X"96",X"16",X"97",X"17",X"0C",X"15",X"26",X"02",X"0C",
		X"14",X"12",X"86",X"14",X"B7",X"20",X"00",X"B6",X"40",X"00",X"C6",X"15",X"F7",X"20",X"01",X"DC",
		X"20",X"2B",X"1F",X"F7",X"60",X"00",X"54",X"4A",X"26",X"13",X"96",X"1F",X"B7",X"78",X"00",X"E6",
		X"A0",X"86",X"08",X"B7",X"78",X"00",X"10",X"9C",X"1D",X"25",X"02",X"86",X"FF",X"DD",X"20",X"F7",
		X"68",X"00",X"DC",X"19",X"3B",X"AA",X"A8",X"54",X"55",X"D5",X"6A",X"55",X"55",X"55",X"B5",X"AA",
		X"20",X"02",X"29",X"A9",X"AD",X"55",X"55",X"95",X"4A",X"55",X"6D",X"DF",X"6D",X"55",X"88",X"90",
		X"A4",X"AA",X"56",X"AB",X"AA",X"AA",X"4A",X"55",X"D5",X"D6",X"EF",X"76",X"55",X"21",X"22",X"51",
		X"AA",X"D6",X"AA",X"AA",X"AA",X"AA",X"52",X"B5",X"BE",X"BB",X"5B",X"55",X"08",X"A1",X"A8",X"AA",
		X"AA",X"55",X"55",X"55",X"55",X"A9",X"6A",X"F3",X"7F",X"AB",X"0A",X"08",X"91",X"AA",X"B5",X"AE",
		X"52",X"A9",X"54",X"A9",X"AA",X"BD",X"EF",X"AE",X"4A",X"00",X"22",X"55",X"DB",X"DA",X"2A",X"A5",
		X"A4",X"54",X"55",X"DF",X"FB",X"5E",X"09",X"01",X"24",X"55",X"F7",X"5A",X"55",X"52",X"92",X"68",
		X"F5",X"7F",X"FF",X"01",X"80",X"D0",X"DF",X"6E",X"40",X"92",X"F6",X"AD",X"12",X"A9",X"FE",X"FF",
		X"03",X"00",X"F8",X"5F",X"2B",X"00",X"AB",X"7F",X"09",X"A2",X"DA",X"FF",X"5D",X"01",X"A0",X"FA",
		X"0F",X"01",X"F8",X"DD",X"26",X"08",X"F6",X"6B",X"77",X"57",X"00",X"58",X"FD",X"A3",X"00",X"BD",
		X"DD",X"09",X"11",X"BE",X"EB",X"ED",X"2D",X"00",X"54",X"FF",X"A1",X"00",X"7D",X"6F",X"41",X"82",
		X"BE",X"DD",X"ED",X"53",X"00",X"58",X"FF",X"21",X"40",X"EF",X"D7",X"20",X"50",X"F7",X"6E",X"7D",
		X"15",X"00",X"D5",X"BF",X"14",X"20",X"B7",X"5F",X"09",X"50",X"DB",X"77",X"FB",X"14",X"00",X"CA",
		X"7F",X"15",X"80",X"B5",X"BF",X"0A",X"90",X"EA",X"EF",X"7E",X"09",X"00",X"EA",X"BF",X"16",X"40",
		X"E5",X"7B",X"2D",X"88",X"A4",X"BF",X"FF",X"14",X"00",X"E4",X"7B",X"2F",X"22",X"A1",X"BA",X"BB",
		X"8A",X"48",X"B5",X"BF",X"2B",X"09",X"90",X"5A",X"5B",X"AD",X"92",X"52",X"AD",X"AA",X"44",X"52",
		X"DB",X"6D",X"AB",X"6A",X"45",X"91",X"AA",X"52",X"A2",X"6A",X"9B",X"A2",X"54",X"7B",X"AB",X"89",
		X"F4",X"AE",X"55",X"B5",X"22",X"91",X"6A",X"AD",X"88",X"A4",X"F6",X"AD",X"22",X"55",X"55",X"55",
		X"7D",X"55",X"44",X"D5",X"AA",X"12",X"29",X"75",X"AD",X"52",X"AA",X"AA",X"4A",X"FB",X"5A",X"85",
		X"AA",X"5A",X"89",X"92",X"DA",X"6A",X"A5",X"AA",X"AA",X"54",X"DD",X"B5",X"A8",X"AA",X"5A",X"89",
		X"22",X"B5",X"AA",X"AA",X"56",X"55",X"52",X"5D",X"55",X"29",X"55",X"5B",X"55",X"11",X"95",X"52",
		X"B5",X"AE",X"48",X"A9",X"AE",X"AA",X"A4",X"AA",X"AE",X"AA",X"92",X"2A",X"AA",X"EA",X"56",X"49",
		X"55",X"AB",X"2A",X"A9",X"AA",X"AE",X"56",X"25",X"95",X"54",X"B5",X"AB",X"4A",X"AA",X"AB",X"52",
		X"A9",X"AA",X"AA",X"AE",X"4A",X"A5",X"94",X"AA",X"AB",X"AA",X"5A",X"55",X"A5",X"AA",X"4A",X"D5",
		X"5B",X"15",X"A5",X"AA",X"6A",X"55",X"A5",X"5A",X"57",X"55",X"51",X"A9",X"AA",X"DF",X"8A",X"A2",
		X"AA",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"29",X"D5",X"AD",X"2A",X"89",X"AA",X"6A",X"55",
		X"55",X"AB",X"AA",X"AA",X"AA",X"A4",X"AA",X"AE",X"AA",X"92",X"AA",X"AA",X"AA",X"AA",X"AB",X"AA",
		X"AA",X"AA",X"52",X"55",X"59",X"55",X"A9",X"2A",X"95",X"AA",X"DA",X"56",X"A9",X"AA",X"55",X"55",
		X"55",X"55",X"D5",X"55",X"AA",X"AA",X"C2",X"B5",X"55",X"47",X"55",X"6A",X"95",X"58",X"AD",X"72",
		X"56",X"13",X"2D",X"4D",X"AE",X"5E",X"A4",X"59",X"4D",X"53",X"A9",X"AA",X"AA",X"AE",X"AA",X"2A",
		X"AA",X"A5",X"74",X"55",X"A3",X"AA",X"9A",X"AA",X"52",X"A5",X"AA",X"AA",X"AA",X"AE",X"F5",X"BD",
		X"BB",X"B7",X"43",X"10",X"14",X"AA",X"EA",X"BA",X"2A",X"89",X"52",X"D5",X"DF",X"FF",X"4A",X"01",
		X"08",X"54",X"F5",X"F5",X"AA",X"22",X"91",X"D4",X"6C",X"F7",X"DD",X"AF",X"18",X"20",X"50",X"D5",
		X"BD",X"5D",X"55",X"50",X"49",X"55",X"AF",X"7B",X"7B",X"4B",X"81",X"10",X"4A",X"ED",X"7A",X"55",
		X"95",X"4A",X"55",X"55",X"55",X"DB",X"B6",X"6D",X"95",X"10",X"49",X"A9",X"52",X"55",X"55",X"55",
		X"AD",X"AA",X"AA",X"EA",X"DE",X"AE",X"55",X"90",X"A4",X"A4",X"28",X"A5",X"AA",X"BA",X"7A",X"B5",
		X"AA",X"5A",X"AF",X"56",X"15",X"89",X"22",X"49",X"94",X"AA",X"6A",X"6D",X"AF",X"56",X"D5",X"54",
		X"55",X"B7",X"2A",X"4A",X"91",X"48",X"92",X"92",X"DA",X"B6",X"B7",X"55",X"29",X"25",X"55",X"75",
		X"BD",X"AD",X"55",X"24",X"49",X"52",X"55",X"AD",X"AA",X"AA",X"AA",X"AA",X"B5",X"BE",X"6B",X"D5",
		X"0A",X"A5",X"52",X"55",X"AD",X"55",X"95",X"12",X"95",X"AA",X"DA",X"56",X"EB",X"C8",X"45",X"55",
		X"AA",X"2A",X"95",X"A2",X"28",X"55",X"A5",X"6A",X"AD",X"D6",X"AA",X"2A",X"29",X"55",X"AA",X"AA",
		X"AA",X"DA",X"AA",X"AA",X"AA",X"AA",X"56",X"55",X"55",X"2A",X"55",X"55",X"55",X"55",X"55",X"55",
		X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"98",X"C3",X"31",X"A3",X"15",X"73",X"1C",
		X"67",X"56",X"8E",X"9C",X"55",X"B9",X"96",X"AA",X"B2",X"94",X"D6",X"54",X"4D",X"73",X"2A",X"A9",
		X"72",X"AC",X"AA",X"19",X"A7",X"2A",X"87",X"8D",X"71",X"C6",X"9C",X"35",X"73",X"CC",X"91",X"39",
		X"4D",X"9A",X"33",X"DB",X"C9",X"A4",X"C6",X"C6",X"19",X"93",X"66",X"C6",X"9C",X"9C",X"33",X"3A",
		X"33",X"E7",X"18",X"6B",X"A6",X"71",X"31",X"B6",X"E1",X"66",X"58",X"8C",X"D9",X"6C",X"8C",X"69",
		X"BB",X"8C",X"2D",X"64",X"5C",X"66",X"CD",X"98",X"63",X"E3",X"2C",X"67",X"C3",X"5C",X"1C",X"67",
		X"F2",X"18",X"8E",X"E3",X"9C",X"99",X"63",X"8E",X"B2",X"34",X"2E",X"E6",X"B2",X"33",X"E7",X"38",
		X"1C",X"C3",X"C8",X"2C",X"6B",X"65",X"96",X"4D",X"D6",X"DD",X"DD",X"99",X"01",X"08",X"93",X"F3",
		X"9D",X"95",X"91",X"92",X"AC",X"7B",X"FF",X"35",X"03",X"02",X"4A",X"5D",X"BF",X"2E",X"09",X"A1",
		X"D4",X"FD",X"FF",X"8A",X"01",X"80",X"AC",X"F7",X"BD",X"14",X"04",X"B1",X"EE",X"FB",X"77",X"20",
		X"00",X"D1",X"F7",X"D7",X"0A",X"08",X"59",X"FD",X"F6",X"6E",X"07",X"04",X"58",X"7F",X"B7",X"08",
		X"48",X"B5",X"77",X"AD",X"EA",X"7E",X"10",X"C0",X"E9",X"BB",X"16",X"08",X"75",X"7D",X"96",X"D4",
		X"F7",X"0F",X"00",X"7C",X"FE",X"49",X"00",X"D9",X"BF",X"09",X"A1",X"FD",X"FF",X"00",X"C0",X"DF",
		X"0F",X"00",X"FC",X"F7",X"02",X"A8",X"FE",X"FB",X"01",X"80",X"FF",X"19",X"00",X"F7",X"1F",X"02",
		X"F1",X"D7",X"DA",X"2E",X"A0",X"E9",X"0F",X"10",X"FA",X"6B",X"01",X"DB",X"B5",X"D0",X"FF",X"03",
		X"28",X"FF",X"80",X"E0",X"3F",X"0A",X"F8",X"93",X"8A",X"FE",X"0F",X"C0",X"FE",X"03",X"E0",X"FE",
		X"80",X"E8",X"2F",X"A8",X"F6",X"3F",X"80",X"7F",X"0F",X"C0",X"7F",X"03",X"78",X"2F",X"A0",X"EF",
		X"3F",X"00",X"FF",X"1C",X"C0",X"DF",X"0A",X"E0",X"5F",X"20",X"FF",X"3F",X"00",X"FE",X"3A",X"00",
		X"FF",X"04",X"E0",X"5F",X"B0",X"FC",X"5F",X"00",X"FF",X"1C",X"80",X"7F",X"41",X"E0",X"1F",X"B4",
		X"F6",X"1F",X"80",X"3F",X"0F",X"C0",X"5F",X"0A",X"F8",X"07",X"B7",X"FD",X"01",X"F0",X"E7",X"00",
		X"F8",X"87",X"06",X"FC",X"A1",X"5F",X"3F",X"00",X"7F",X"1C",X"80",X"FF",X"A0",X"C0",X"9F",X"E8",
		X"BF",X"02",X"F0",X"4F",X"02",X"F8",X"0F",X"09",X"FA",X"95",X"FE",X"0B",X"80",X"7F",X"25",X"C0",
		X"7F",X"09",X"C1",X"7E",X"B5",X"3F",X"00",X"FE",X"69",X"00",X"FE",X"53",X"04",X"FA",X"5B",X"FF",
		X"00",X"F8",X"A7",X"05",X"F0",X"4F",X"1A",X"E0",X"3F",X"FD",X"01",X"F0",X"4F",X"0B",X"C0",X"7F",
		X"38",X"00",X"FF",X"EB",X"03",X"E0",X"1F",X"1E",X"80",X"FF",X"A8",X"04",X"FE",X"5F",X"01",X"E0",
		X"7F",X"14",X"00",X"FF",X"13",X"81",X"FE",X"7F",X"00",X"F0",X"BF",X"11",X"80",X"FF",X"95",X"00",
		X"FF",X"1F",X"00",X"FE",X"76",X"01",X"E8",X"75",X"97",X"A0",X"FF",X"00",X"A8",X"FB",X"2B",X"00",
		X"7D",X"57",X"A5",X"F6",X"03",X"B0",X"CB",X"BD",X"80",X"54",X"F5",X"2D",X"FD",X"05",X"80",X"B7",
		X"DD",X"02",X"52",X"6B",X"55",X"FF",X"0F",X"00",X"DC",X"7B",X"05",X"52",X"D5",X"6A",X"FB",X"3F",
		X"00",X"58",X"FB",X"0B",X"50",X"B2",X"5D",X"FB",X"3F",X"00",X"54",X"FE",X"05",X"95",X"50",X"DB",
		X"FF",X"17",X"00",X"AA",X"BF",X"A0",X"45",X"D8",X"B6",X"FB",X"07",X"00",X"EA",X"BF",X"88",X"90",
		X"DA",X"EE",X"BF",X"00",X"20",X"F5",X"5B",X"4B",X"80",X"DA",X"FF",X"0F",X"00",X"CA",X"6D",X"B5",
		X"0A",X"45",X"F5",X"FF",X"45",X"00",X"D8",X"DD",X"26",X"52",X"52",X"EF",X"3F",X"11",X"88",X"AA",
		X"B6",X"25",X"25",X"A9",X"BF",X"AF",X"08",X"91",X"B4",X"76",X"05",X"A5",X"BA",X"76",X"AB",X"CA",
		X"44",X"61",X"66",X"33",X"41",X"AB",X"7A",X"B5",X"AA",X"91",X"5E",X"16",X"89",X"B5",X"AA",X"88",
		X"A6",X"55",X"35",X"4B",X"57",X"12",X"31",X"2D",X"95",X"2A",X"55",X"B5",X"AA",X"9A",X"64",X"92",
		X"A6",X"B8",X"2C",X"45",X"D6",X"B6",X"A8",X"9A",X"62",X"BA",X"54",X"95",X"44",X"D7",X"AA",X"52",
		X"A5",X"6A",X"35",X"6B",X"11",X"52",X"B5",X"AB",X"52",X"55",X"51",X"A9",X"6A",X"A9",X"AA",X"B5",
		X"DA",X"A8",X"50",X"4B",X"D3",X"A8",X"26",X"95",X"DA",X"AD",X"50",X"29",X"6B",X"15",X"A5",X"AA",
		X"B5",X"2A",X"65",X"A5",X"6A",X"55",X"A5",X"AA",X"AA",X"66",X"B6",X"52",X"4B",X"55",X"2D",X"6A",
		X"A7",X"CA",X"52",X"45",X"55",X"B6",X"55",X"A2",X"6A",X"5D",X"2A",X"99",X"AD",X"05",X"AD",X"74",
		X"53",X"58",X"CB",X"CA",X"95",X"AA",X"AA",X"56",X"D3",X"5A",X"55",X"49",X"AB",X"93",X"52",X"5B",
		X"AA",X"2D",X"A9",X"F6",X"2A",X"55",X"95",X"22",X"55",X"6D",X"A9",X"2A",X"AD",X"DA",X"32",X"15",
		X"B6",X"2A",X"5D",X"4A",X"59",X"35",X"5D",X"4B",X"A9",X"54",X"D5",X"EA",X"52",X"29",X"AB",X"6A",
		X"69",X"49",X"B2",X"6A",X"D5",X"AC",X"68",X"5B",X"B2",X"6A",X"54",X"B4",X"CA",X"55",X"5A",X"51",
		X"D5",X"6C",X"55",X"AA",X"54",X"D5",X"AA",X"A9",X"E4",X"AA",X"D2",X"75",X"AB",X"54",X"55",X"AA",
		X"56",X"25",X"55",X"A5",X"5A",X"95",X"AA",X"74",X"D5",X"56",X"A2",X"C5",X"AA",X"95",X"95",X"46",
		X"4B",X"AA",X"5E",X"55",X"59",X"B5",X"54",X"51",X"55",X"AB",X"BA",X"52",X"29",X"B5",X"4A",X"52",
		X"6B",X"AD",X"94",X"5C",X"AB",X"34",X"55",X"A9",X"AA",X"CB",X"B6",X"AA",X"4A",X"55",X"52",X"55",
		X"55",X"55",X"AD",X"B5",X"AC",X"DC",X"AA",X"4A",X"55",X"AA",X"A5",X"55",X"55",X"B4",X"A4",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"56",X"2D",X"55",X"55",X"55",X"55",X"53",X"A4",X"A6",
		X"AA",X"B5",X"B2",X"56",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"6A",X"2B",X"15",X"A9",X"E9",X"AA",X"AA",X"D6",X"2A",X"A9",X"AA",X"54",X"55",
		X"55",X"B5",X"5A",X"55",X"55",X"4A",X"AB",X"AA",X"5A",X"55",X"95",X"AA",X"AA",X"AA",X"AA",X"5A",
		X"55",X"55",X"65",X"55",X"A5",X"A6",X"AA",X"6D",X"29",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"52",X"55",X"55",X"AB",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AD",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"52",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AB",
		X"AA",X"4C",X"B6",X"6C",X"9C",X"2E",X"55",X"D9",X"64",X"CE",X"8E",X"C1",X"CC",X"66",X"B7",X"91",
		X"26",X"4B",X"A6",X"6A",X"B2",X"36",X"AD",X"55",X"B2",X"34",X"D3",X"28",X"D9",X"94",X"66",X"ED",
		X"DA",X"B6",X"6D",X"12",X"48",X"92",X"C3",X"72",X"B3",X"9F",X"9F",X"CD",X"08",X"44",X"CC",X"AA",
		X"95",X"35",X"EF",X"7D",X"3D",X"0A",X"84",X"D0",X"74",X"BD",X"55",X"65",X"DD",X"D7",X"C5",X"40",
		X"40",X"CA",X"EB",X"5B",X"0B",X"D7",X"3E",X"0F",X"07",X"04",X"2A",X"AF",X"AF",X"56",X"AA",X"7B",
		X"7C",X"0C",X"10",X"68",X"7C",X"5F",X"73",X"54",X"FE",X"38",X"3C",X"40",X"C8",X"BC",X"BE",X"5A",
		X"94",X"FE",X"F0",X"38",X"08",X"B0",X"F8",X"7C",X"AD",X"18",X"BD",X"E3",X"71",X"10",X"50",X"E5",
		X"FD",X"5C",X"94",X"F4",X"8F",X"E3",X"41",X"40",X"AA",X"FB",X"B5",X"A4",X"E8",X"3D",X"1E",X"07",
		X"01",X"A9",X"D7",X"AF",X"89",X"A2",X"7F",X"3C",X"0E",X"04",X"94",X"5E",X"5F",X"47",X"8A",X"FE",
		X"F1",X"38",X"10",X"50",X"6E",X"DF",X"9A",X"12",X"ED",X"C7",X"E3",X"20",X"20",X"D9",X"7D",X"AB",
		X"A2",X"F4",X"1E",X"8F",X"83",X"80",X"E2",X"F6",X"AE",X"8A",X"B2",X"3F",X"1E",X"07",X"01",X"C5",
		X"EE",X"6D",X"53",X"E4",X"FE",X"78",X"1C",X"04",X"84",X"DB",X"B7",X"A6",X"94",X"FD",X"F1",X"38",
		X"08",X"28",X"3B",X"9F",X"8B",X"51",X"F7",X"E7",X"A1",X"20",X"30",X"DD",X"9E",X"16",X"C6",X"F6",
		X"3F",X"07",X"81",X"A0",X"B5",X"75",X"55",X"68",X"BC",X"FF",X"39",X"08",X"04",X"AB",X"D3",X"69",
		X"52",X"DA",X"FD",X"CF",X"01",X"30",X"58",X"AE",X"56",X"25",X"D5",X"EE",X"BF",X"07",X"40",X"B0",
		X"6A",X"B5",X"96",X"94",X"F5",X"FF",X"1C",X"04",X"82",X"A5",X"B3",X"B5",X"A4",X"EA",X"FF",X"F3",
		X"00",X"08",X"96",X"55",X"D7",X"A2",X"B4",X"FE",X"CF",X"43",X"20",X"A8",X"9C",X"AD",X"A5",X"A4",
		X"FD",X"3F",X"0F",X"80",X"41",X"B5",X"6A",X"4B",X"A9",X"EA",X"FF",X"3C",X"04",X"82",X"CA",X"AA",
		X"AB",X"52",X"DA",X"FF",X"E7",X"20",X"08",X"4A",X"AB",X"5A",X"8D",X"AA",X"FE",X"9F",X"43",X"20",
		X"28",X"AD",X"5A",X"A7",X"E2",X"FC",X"3F",X"07",X"41",X"21",X"6A",X"B5",X"56",X"C6",X"EA",X"FF",
		X"3C",X"04",X"82",X"58",X"55",X"AB",X"2A",X"AB",X"FF",X"73",X"28",X"08",X"92",X"55",X"6B",X"A5",
		X"AC",X"FE",X"EF",X"41",X"20",X"28",X"55",X"AD",X"95",X"A9",X"FE",X"3F",X"87",X"40",X"50",X"AC",
		X"6A",X"2D",X"47",X"F3",X"FF",X"1C",X"0A",X"82",X"64",X"55",X"AD",X"2A",X"AB",X"FF",X"73",X"18",
		X"08",X"A1",X"59",X"D5",X"AA",X"AA",X"FE",X"CF",X"61",X"20",X"88",X"A6",X"6A",X"AB",X"AA",X"F5",
		X"BF",X"46",X"81",X"20",X"1C",X"AB",X"56",X"55",X"ED",X"F7",X"1D",X"0A",X"82",X"D0",X"54",X"6D",
		X"55",X"56",X"FF",X"D7",X"28",X"08",X"42",X"A5",X"EA",X"6A",X"59",X"7D",X"BF",X"47",X"41",X"10",
		X"1C",X"AB",X"D5",X"AA",X"B9",X"F7",X"5D",X"04",X"81",X"E0",X"58",X"AD",X"56",X"55",X"EF",X"EF",
		X"28",X"08",X"84",X"A6",X"6A",X"AD",X"AA",X"EE",X"EF",X"A6",X"40",X"10",X"54",X"56",X"57",X"55",
		X"B5",X"DF",X"B7",X"04",X"02",X"A1",X"52",X"5D",X"97",X"6A",X"FB",X"BE",X"55",X"20",X"10",X"4A",
		X"CB",X"B5",X"AA",X"76",X"FF",X"2E",X"05",X"81",X"50",X"AA",X"AE",X"55",X"D5",X"FD",X"DE",X"8A",
		X"10",X"80",X"52",X"B5",X"B5",X"AA",X"F6",X"FB",X"56",X"41",X"00",X"49",X"5A",X"AB",X"55",X"6D",
		X"BF",X"6F",X"25",X"10",X"20",X"A9",X"DA",X"5A",X"D5",X"F6",X"DF",X"55",X"02",X"02",X"92",X"AA",
		X"AD",X"AB",X"DA",X"FB",X"5B",X"45",X"00",X"90",X"AA",X"5A",X"5B",X"AD",X"FB",X"B7",X"95",X"00",
		X"40",X"52",X"B5",X"B6",X"EA",X"7A",X"7F",X"5B",X"02",X"02",X"A4",X"AA",X"B6",X"AD",X"D6",X"FB",
		X"D7",X"12",X"08",X"20",X"55",X"75",X"5D",X"AD",X"7D",X"DF",X"2A",X"02",X"80",X"94",X"6A",X"EB",
		X"6A",X"ED",X"DF",X"56",X"11",X"00",X"24",X"D5",X"DA",X"6A",X"6D",X"FF",X"6D",X"29",X"00",X"84",
		X"52",X"6B",X"AB",X"B5",X"FD",X"B7",X"95",X"40",X"00",X"2A",X"AD",X"6D",X"AD",X"F6",X"FD",X"36",
		X"0A",X"00",X"A2",X"AA",X"DA",X"56",X"EB",X"FE",X"6D",X"45",X"00",X"84",X"54",X"AD",X"AD",X"D5",
		X"EE",X"DF",X"2A",X"01",X"20",X"54",X"5A",X"5B",X"5B",X"DB",X"7F",X"5B",X"12",X"00",X"24",X"55",
		X"6B",X"AB",X"6D",X"FF",X"DB",X"92",X"00",X"20",X"A9",X"6A",X"6D",X"AD",X"7D",X"7F",X"2B",X"01",
		X"01",X"92",X"AA",X"B5",X"56",X"BB",X"FF",X"B6",X"24",X"00",X"48",X"AA",X"DA",X"5A",X"6B",X"DF",
		X"DF",X"4A",X"04",X"40",X"54",X"D5",X"5A",X"5B",X"FB",X"DF",X"2E",X"09",X"00",X"92",X"AA",X"D6",
		X"6A",X"DB",X"FE",X"DB",X"12",X"01",X"20",X"AA",X"AA",X"AD",X"D6",X"EE",X"DF",X"96",X"04",X"00",
		X"49",X"55",X"6B",X"75",X"ED",X"FE",X"6D",X"09",X"08",X"08",X"55",X"B5",X"56",X"DB",X"EE",X"DF",
		X"A6",X"00",X"20",X"52",X"55",X"6B",X"B5",X"DD",X"BF",X"5B",X"12",X"00",X"22",X"55",X"6D",X"B5",
		X"B5",X"FB",X"B7",X"25",X"01",X"40",X"54",X"55",X"5B",X"5B",X"7B",X"7F",X"57",X"02",X"02",X"44",
		X"D5",X"6A",X"AD",X"6D",X"FF",X"6D",X"25",X"40",X"40",X"AA",X"6A",X"AD",X"B6",X"7D",X"BF",X"2D",
		X"02",X"80",X"A4",X"AA",X"B6",X"D6",X"B6",X"FF",X"B6",X"24",X"00",X"88",X"AA",X"5A",X"AB",X"6D",
		X"FB",X"6F",X"4B",X"02",X"80",X"A8",X"AA",X"AD",X"B6",X"76",X"FF",X"B6",X"24",X"00",X"48",X"AA",
		X"D6",X"5A",X"6D",X"F7",X"6F",X"4B",X"02",X"80",X"A8",X"6A",X"AD",X"AE",X"B6",X"BF",X"5B",X"09",
		X"00",X"44",X"AA",X"B5",X"D5",X"DA",X"EE",X"6F",X"2B",X"01",X"80",X"A8",X"6A",X"6D",X"AB",X"6D",
		X"FF",X"B6",X"12",X"00",X"88",X"AA",X"D6",X"D6",X"5A",X"FB",X"BE",X"2D",X"01",X"80",X"C8",X"AA",
		X"B5",X"6D",X"6D",X"EF",X"DB",X"8A",X"00",X"40",X"AA",X"6A",X"DB",X"D6",X"B6",X"DF",X"B5",X"04",
		X"08",X"A0",X"AA",X"DA",X"B6",X"B5",X"DD",X"B7",X"96",X"02",X"20",X"A4",X"AA",X"B6",X"5D",X"5B",
		X"F7",X"56",X"55",X"21",X"20",X"52",X"AA",X"B6",X"6E",X"6B",X"6B",X"AB",X"55",X"15",X"04",X"91",
		X"A4",X"6A",X"DB",X"6D",X"AB",X"B5",X"D6",X"AA",X"42",X"20",X"24",X"55",X"B5",X"75",X"AD",X"56",
		X"B5",X"DD",X"AE",X"0A",X"42",X"48",X"2A",X"B5",X"6A",X"5D",X"95",X"AA",X"BB",X"AE",X"55",X"41",
		X"28",X"52",X"AA",X"AA",X"AA",X"AA",X"AA",X"BD",X"BB",X"AD",X"0A",X"91",X"48",X"4A",X"A5",X"AA",
		X"6A",X"ED",X"D5",X"DA",X"5A",X"AB",X"42",X"92",X"28",X"A5",X"AA",X"AA",X"5A",X"55",X"55",X"55",
		X"AD",X"6F",X"AB",X"22",X"8A",X"44",X"4A",X"AA",X"AA",X"D6",X"AA",X"AA",X"AA",X"EA",X"BB",X"AA",
		X"10",X"51",X"52",X"55",X"55",X"55",X"55",X"5D",X"55",X"55",X"52",X"55",X"D5",X"6A",X"55",X"8A",
		X"92",X"52",X"52",X"AA",X"6A",X"AB",X"5A",X"55",X"55",X"55",X"2A",X"8A",X"52",X"52",X"D5",X"D6",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"4A",X"55",X"55",X"55",X"55",X"55",X"B5",X"AA",X"AA",
		X"A4",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"D5",
		X"AA",X"94",X"AA",X"E2",X"55",X"5D",X"A5",X"AA",X"2A",X"55",X"55",X"A9",X"54",X"11",X"2E",X"FD",
		X"BB",X"4A",X"A3",X"AA",X"7A",X"EB",X"BA",X"55",X"15",X"22",X"A1",X"54",X"AD",X"6F",X"77",X"F7",
		X"17",X"07",X"02",X"20",X"6A",X"F5",X"DD",X"14",X"45",X"B5",X"FF",X"7C",X"18",X"40",X"20",X"AB",
		X"F7",X"B5",X"95",X"A4",X"EE",X"CB",X"E3",X"81",X"80",X"A8",X"AE",X"9F",X"97",X"C3",X"72",X"2F",
		X"1F",X"07",X"06",X"C2",X"BA",X"BE",X"9E",X"26",X"A6",X"BD",X"7C",X"1C",X"0C",X"04",X"CE",X"BE",
		X"3B",X"17",X"0D",X"D7",X"E5",X"71",X"30",X"10",X"1C",X"7B",X"BB",X"AD",X"4A",X"6A",X"0F",X"8F",
		X"87",X"81",X"C0",X"E9",X"F5",X"75",X"69",X"D2",X"7C",X"78",X"1C",X"0C",X"12",X"0E",X"AF",X"D7",
		X"55",X"45",X"F5",X"C5",X"E3",X"60",X"10",X"B1",X"78",X"BE",X"9E",X"96",X"54",X"6F",X"3C",X"0E",
		X"06",X"09",X"D3",X"D3",X"FB",X"B8",X"64",X"7A",X"D5",X"E3",X"50",X"10",X"38",X"7A",X"BE",X"AB",
		X"25",X"A5",X"D7",X"3C",X"0E",X"03",X"81",X"A9",X"E7",X"DB",X"5A",X"32",X"7A",X"CB",X"E3",X"50",
		X"10",X"98",X"BA",X"BE",X"AE",X"A5",X"C6",X"6D",X"3D",X"0E",X"06",X"81",X"C5",X"F3",X"75",X"B5",
		X"2A",X"DA",X"2D",X"C7",X"E1",X"20",X"30",X"DA",X"7A",X"2F",X"A7",X"CA",X"DA",X"F1",X"38",X"1C",
		X"04",X"26",X"97",X"D7",X"F3",X"68",X"AC",X"AE",X"3C",X"0E",X"07",X"A1",X"62",X"F5",X"DC",X"5A",
		X"55",X"D5",X"56",X"8F",X"C3",X"41",X"50",X"B4",X"3C",X"AF",X"96",X"D5",X"72",X"35",X"CF",X"C5",
		X"20",X"28",X"AC",X"5A",X"AB",X"4E",X"AB",X"71",X"75",X"BA",X"2E",X"83",X"20",X"51",X"D5",X"6A",
		X"39",X"2D",X"AD",X"D6",X"F5",X"E9",X"32",X"28",X"28",X"55",X"4D",X"4B",X"55",X"55",X"5D",X"AF",
		X"ED",X"5A",X"15",X"8A",X"A2",X"4A",X"A5",X"A8",X"54",X"ED",X"75",X"AD",X"DA",X"76",X"AD",X"14",
		X"0A",X"85",X"44",X"AA",X"6A",X"EB",X"AA",X"AA",X"EA",X"BB",X"5B",X"15",X"44",X"48",X"4A",X"55",
		X"55",X"B5",X"5A",X"75",X"DB",X"DE",X"B6",X"2A",X"41",X"92",X"94",X"52",X"52",X"AA",X"B6",X"6F",
		X"6B",X"55",X"AD",X"6B",X"B5",X"10",X"12",X"29",X"25",X"55",X"D5",X"B6",X"BA",X"4A",X"55",X"F5",
		X"BA",X"56",X"21",X"89",X"94",X"52",X"A9",X"AA",X"AA",X"AD",X"AA",X"AA",X"AA",X"AA",X"7A",X"AD",
		X"88",X"A2",X"A8",X"94",X"52",X"55",X"AD",X"DD",X"AA",X"52",X"2A",X"55",X"D5",X"DA",X"AA",X"8A",
		X"52",X"55",X"55",X"A5",X"52",X"A9",X"AA",X"55",X"55",X"55",X"55",X"B5",X"75",X"7D",X"AB",X"A5",
		X"4A",X"8A",X"92",X"28",X"A9",X"AA",X"B6",X"B5",X"AA",X"AA",X"77",X"5D",X"AB",X"42",X"22",X"92",
		X"4A",X"55",X"E1",X"3C",X"7A",X"AD",X"56",X"B9",X"4A",X"A5",X"38",X"96",X"8A",X"E3",X"78",X"C4",
		X"39",X"CE",X"E5",X"1C",X"C7",X"11",X"A7",X"73",X"9C",X"71",X"28",X"96",X"29",X"E7",X"56",X"C5",
		X"99",X"9A",X"B7",X"B6",X"2A",X"24",X"8A",X"52",X"55",X"AD",X"AB",X"39",X"C6",X"AA",X"BB",X"F3",
		X"2C",X"10",X"24",X"4C",X"6D",X"AF",X"AD",X"2A",X"A5",X"F6",X"B7",X"9E",X"03",X"02",X"A1",X"AA",
		X"EB",X"DB",X"AA",X"A2",X"EE",X"3B",X"C7",X"81",X"80",X"C4",X"F4",X"DE",X"6B",X"A9",X"A8",X"FE",
		X"F2",X"1C",X"10",X"50",X"8C",X"7B",X"5F",X"8D",X"28",X"F5",X"8F",X"C7",X"01",X"01",X"C3",X"ED",
		X"7B",X"55",X"42",X"B1",X"7F",X"79",X"06",X"08",X"18",X"BE",X"7E",X"4F",X"0A",X"8A",X"FD",X"D7",
		X"63",X"00",X"C0",X"F1",X"FB",X"AD",X"21",X"50",X"FA",X"3F",X"1E",X"03",X"00",X"CD",X"DF",X"AF",
		X"0A",X"02",X"EB",X"FF",X"EB",X"00",X"80",X"F0",X"FA",X"7B",X"45",X"20",X"B8",X"FD",X"7F",X"1C",
		X"00",X"48",X"BD",X"7F",X"87",X"00",X"4A",X"FF",X"FF",X"0B",X"03",X"80",X"D5",X"EF",X"D3",X"00",
		X"A1",X"EB",X"FB",X"B7",X"60",X"00",X"BC",X"F5",X"74",X"18",X"6A",X"5C",X"BA",X"FE",X"3D",X"0C",
		X"80",X"B6",X"1E",X"1D",X"8B",X"96",X"2C",X"B6",X"FE",X"3F",X"0C",X"00",X"BB",X"1E",X"1F",X"0A",
		X"17",X"2D",X"5D",X"FF",X"1F",X"04",X"80",X"B7",X"1E",X"17",X"1C",X"1D",X"56",X"5D",X"7F",X"1F",
		X"0C",X"00",X"7F",X"1E",X"19",X"35",X"35",X"59",X"5A",X"FF",X"7D",X"30",X"00",X"FE",X"74",X"A8",
		X"D4",X"E2",X"A8",X"AA",X"F7",X"BF",X"81",X"80",X"F8",X"C7",X"C1",X"A2",X"95",X"C3",X"B1",X"AD",
		X"DF",X"0F",X"04",X"4C",X"3F",X"1C",X"AC",X"3C",X"5C",X"B8",X"BC",X"FA",X"BE",X"42",X"60",X"FA",
		X"C3",X"60",X"95",X"47",X"25",X"AB",X"AE",X"F7",X"3B",X"08",X"4C",X"77",X"18",X"8C",X"F3",X"A8",
		X"D1",X"D4",X"E9",X"FB",X"0B",X"03",X"CB",X"1D",X"02",X"67",X"5D",X"95",X"A2",X"AA",X"EE",X"FF",
		X"07",X"81",X"4A",X"0F",X"83",X"6B",X"5D",X"8A",X"C2",X"DA",X"DD",X"BF",X"07",X"02",X"4E",X"1F",
		X"0A",X"67",X"35",X"52",X"B2",X"76",X"AB",X"F7",X"1F",X"04",X"6C",X"7C",X"48",X"78",X"79",X"A8",
		X"98",X"D6",X"5A",X"7E",X"FF",X"20",X"60",X"E3",X"43",X"45",X"8F",X"16",X"4E",X"1E",X"5D",X"B9",
		X"FE",X"0E",X"04",X"6E",X"3C",X"94",X"E4",X"B1",X"45",X"47",X"8D",X"55",X"BD",X"FF",X"05",X"80",
		X"1B",X"0F",X"15",X"75",X"3C",X"52",X"71",X"55",X"A7",X"EB",X"BE",X"05",X"C0",X"36",X"1E",X"52",
		X"78",X"75",X"52",X"69",X"A9",X"55",X"D7",X"FD",X"07",X"00",X"3B",X"1E",X"52",X"E9",X"A9",X"91",
		X"A6",X"36",X"1E",X"55",X"FD",X"3B",X"00",X"F8",X"E3",X"20",X"15",X"5F",X"2D",X"34",X"E5",X"64",
		X"A5",X"EB",X"7E",X"07",X"00",X"3F",X"1E",X"52",X"E5",X"A5",X"86",X"66",X"2D",X"96",X"B4",X"FA",
		X"B7",X"03",X"80",X"1F",X"1E",X"B2",X"F8",X"4A",X"C1",X"AA",X"2D",X"2A",X"B5",X"F9",X"6D",X"07",
		X"84",X"7E",X"58",X"D0",X"D1",X"8B",X"8A",X"5A",X"75",X"A8",X"AA",X"CB",X"DB",X"3E",X"20",X"E8",
		X"A5",X"06",X"55",X"5A",X"55",X"A9",X"56",X"17",X"4A",X"5A",X"F5",X"F7",X"0D",X"90",X"B8",X"A2",
		X"92",X"1A",X"BD",X"68",X"A9",X"4B",X"45",X"6A",X"76",X"D5",X"D7",X"AF",X"20",X"48",X"55",X"5A",
		X"D2",X"AA",X"55",X"95",X"AA",X"4A",X"59",X"55",X"4D",X"DD",X"EE",X"5E",X"55",X"41",X"90",X"A8",
		X"54",X"55",X"55",X"B5",X"AE",X"4A",X"55",X"A4",X"64",X"D7",X"DF",X"5E",X"29",X"10",X"44",X"4A",
		X"55",X"D5",X"AA",X"BA",X"AD",X"2A",X"29",X"4A",X"55",X"F7",X"DE",X"B6",X"84",X"10",X"22",X"A9",
		X"AA",X"F5",X"AA",X"5A",X"AB",X"54",X"54",X"AA",X"AA",X"DD",X"DB",X"AD",X"04",X"09",X"A2",X"A4",
		X"AA",X"5A",X"AD",X"AA",X"AA",X"4A",X"25",X"A5",X"6A",X"FD",X"EE",X"B6",X"0A",X"21",X"24",X"A9",
		X"54",X"B5",X"5A",X"DD",X"5A",X"55",X"4A",X"55",X"AA",X"FA",X"ED",X"B5",X"2A",X"24",X"88",X"A8",
		X"AA",X"AA",X"5A",X"BB",X"B6",X"AA",X"22",X"55",X"55",X"B5",X"F7",X"B6",X"2A",X"88",X"48",X"94",
		X"AA",X"AA",X"5A",X"AD",X"AA",X"AA",X"54",X"AA",X"AA",X"DA",X"BE",X"AE",X"AB",X"82",X"10",X"49",
		X"A9",X"52",X"B5",X"6A",X"75",X"A9",X"AA",X"52",X"2A",X"D5",X"BE",X"BB",X"AD",X"12",X"82",X"90",
		X"54",X"55",X"AD",X"6A",X"55",X"55",X"55",X"55",X"AA",X"6A",X"EF",X"ED",X"5A",X"05",X"21",X"91",
		X"54",X"55",X"D5",X"6A",X"55",X"57",X"B5",X"54",X"95",X"AA",X"F6",X"DD",X"56",X"85",X"10",X"89",
		X"A4",X"AA",X"AA",X"D5",X"AA",X"6B",X"55",X"AA",X"AA",X"AA",X"BE",X"DE",X"5A",X"15",X"44",X"42",
		X"49",X"55",X"D5",X"5A",X"55",X"75",X"AD",X"4A",X"55",X"B5",X"DB",X"F6",X"6A",X"15",X"44",X"44",
		X"94",X"AA",X"AA",X"6A",X"B5",X"AA",X"52",X"55",X"55",X"55",X"ED",X"DD",X"56",X"15",X"22",X"42",
		X"92",X"4A",X"55",X"AB",X"55",X"57",X"A9",X"AA",X"AA",X"EA",X"75",X"5D",X"5B",X"AB",X"90",X"08",
		X"49",X"AA",X"AA",X"5A",X"AB",X"53",X"55",X"55",X"95",X"6A",X"F5",X"AE",X"6D",X"B5",X"0A",X"09",
		X"91",X"A8",X"AA",X"AA",X"5A",X"AD",X"AA",X"AA",X"AA",X"AA",X"BA",X"DB",X"76",X"5B",X"55",X"21",
		X"22",X"4A",X"A9",X"AA",X"5A",X"55",X"AB",X"AA",X"AA",X"AA",X"AA",X"DE",X"AE",X"5B",X"AB",X"42",
		X"22",X"92",X"A4",X"54",X"55",X"55",X"AB",X"AA",X"AA",X"AA",X"52",X"55",X"5B",X"AB",X"B7",X"92",
		X"88",X"84",X"A4",X"54",X"AA",X"AA",X"6A",X"B5",X"AA",X"AA",X"AA",X"AA",X"56",X"BF",X"6D",X"5B",
		X"55",X"91",X"24",X"92",X"52",X"A9",X"AA",X"AE",X"AA",X"AA",X"AA",X"AA",X"AA",X"F5",X"6E",X"D7",
		X"AA",X"2A",X"8A",X"22",X"51",X"AA",X"54",X"55",X"AB",X"56",X"55",X"55",X"55",X"AD",X"DE",X"D6",
		X"6A",X"29",X"8A",X"A2",X"A8",X"A8",X"AA",X"AA",X"6A",X"55",X"55",X"55",X"55",X"B5",X"D6",X"B7",
		X"B6",X"5A",X"2D",X"52",X"92",X"24",X"4A",X"A5",X"AA",X"AA",X"56",X"55",X"55",X"55",X"6B",X"B5",
		X"5A",X"55",X"49",X"92",X"24",X"44",X"52",X"52",X"55",X"AD",X"5A",X"B5",X"AA",X"AA",X"AA",X"B6",
		X"AA",X"AA",X"77",X"29",X"95",X"52",X"49",X"55",X"D5",X"EA",X"6A",X"55",X"0F",X"FB",X"A1",X"6A",
		X"F4",X"6A",X"95",X"2A",X"95",X"2B",X"55",X"7A",X"A5",X"DA",X"6A",X"2D",X"B5",X"56",X"5A",X"69",
		X"B5",X"94",X"50",X"42",X"A9",X"94",X"56",X"6B",X"A5",X"D5",X"EA",X"F5",X"EB",X"E1",X"C0",X"A0",
		X"50",X"D5",X"6A",X"A7",X"43",X"A3",X"12",X"A5",X"56",X"AF",X"D7",X"6B",X"97",X"16",X"05",X"85",
		X"96",X"5A",X"6B",X"BD",X"96",X"12",X"6A",X"38",X"3D",X"B7",X"7B",X"AF",X"D6",X"A0",X"50",X"28",
		X"D5",X"EA",X"DD",X"5A",X"15",X"4A",X"38",X"16",X"AF",X"D7",X"6B",X"AF",X"16",X"05",X"85",X"44",
		X"56",X"6B",X"AF",X"A5",X"94",X"42",X"C2",X"71",X"B5",X"FD",X"7A",X"3D",X"0E",X"0A",X"41",X"A9",
		X"9C",X"EB",X"E5",X"52",X"A1",X"50",X"2A",X"9D",X"DE",X"6B",X"AF",X"E5",X"30",X"08",X"0A",X"2B",
		X"BD",X"9E",X"97",X"4A",X"0A",X"25",X"A5",X"F3",X"76",X"EF",X"D6",X"3A",X"04",X"0A",X"A5",X"4A",
		X"AF",X"D7",X"AA",X"14",X"29",X"94",X"4E",X"AF",X"77",X"AF",X"D7",X"60",X"21",X"18",X"6A",X"79",
		X"3D",X"3D",X"55",X"92",X"42",X"4B",X"ED",X"F5",X"F6",X"7A",X"55",X"18",X"04",X"16",X"AB",X"56",
		X"AF",X"C7",X"62",X"28",X"4A",X"65",X"F5",X"6E",X"AF",X"B5",X"0A",X"81",X"C1",X"D0",X"D2",X"DA",
		X"79",X"29",X"25",X"94",X"92",X"D6",X"5E",X"EF",X"AD",X"56",X"0A",X"04",X"49",X"A5",X"D6",X"EB",
		X"56",X"23",X"25",X"52",X"A5",X"D5",X"6F",X"EF",X"D5",X"52",X"01",X"A1",X"C4",X"F2",X"F2",X"5A",
		X"4B",X"29",X"29",X"A5",X"B4",X"F5",X"DE",X"7B",X"B5",X"18",X"08",X"94",X"4A",X"AD",X"75",X"AB",
		X"A5",X"14",X"29",X"95",X"56",X"DF",X"ED",X"D7",X"4A",X"09",X"84",X"A4",X"D4",X"D6",X"D6",X"4B",
		X"4B",X"28",X"29",X"AD",X"BC",X"BD",X"DE",X"4B",X"C7",X"40",X"28",X"D1",X"58",X"AD",X"75",X"5A",
		X"25",X"12",X"4B",X"A5",X"F5",X"5E",X"6F",X"AD",X"D1",X"20",X"18",X"4A",X"5A",X"5B",X"2F",X"2D",
		X"25",X"A5",X"A4",X"A5",X"F5",X"BD",X"5E",X"6B",X"34",X"08",X"0A",X"A5",X"5A",X"8F",X"D7",X"52",
		X"29",X"52",X"4A",X"B3",X"F5",X"7A",X"AF",X"35",X"1A",X"02",X"61",X"A9",X"B5",X"B5",X"B5",X"96",
		X"42",X"52",X"6A",X"5A",X"7B",X"AF",X"B7",X"5A",X"0C",X"06",X"42",X"A5",X"D5",X"6B",X"B5",X"52",
		X"2A",X"85",X"CA",X"69",X"BD",X"D7",X"5E",X"2D",X"06",X"42",X"22",X"AB",X"B5",X"7A",X"5A",X"A5",
		X"14",X"4A",X"A5",X"D5",X"BB",X"D7",X"55",X"A3",X"A0",X"10",X"55",X"5C",X"55",X"D7",X"A9",X"A8",
		X"A8",X"AA",X"AA",X"BE",X"5D",X"57",X"1D",X"83",X"A1",X"28",X"56",X"ED",X"5A",X"95",X"A3",X"68",
		X"94",X"AA",X"57",X"AF",X"EB",X"AA",X"08",X"85",X"44",X"55",X"D5",X"75",X"B5",X"8A",X"AA",X"A8",
		X"AA",X"56",X"5F",X"DF",X"E5",X"28",X"08",X"45",X"AA",X"56",X"E7",X"6A",X"55",X"2A",X"52",X"C5",
		X"AA",X"77",X"7D",X"B5",X"AA",X"20",X"28",X"46",X"6B",X"55",X"75",X"55",X"2C",X"2A",X"AA",X"EA",
		X"D5",X"F5",X"B5",X"AA",X"42",X"41",X"A9",X"2A",X"75",X"AD",X"4B",X"B5",X"28",X"55",X"A9",X"DA",
		X"F5",X"75",X"B5",X"38",X"28",X"8A",X"A2",X"E5",X"71",X"75",X"55",X"54",X"45",X"D5",X"AA",X"EA",
		X"AE",X"57",X"55",X"85",X"A2",X"54",X"B4",X"AA",X"55",X"AB",X"4A",X"55",X"AA",X"6A",X"55",X"BD",
		X"AA",X"AB",X"63",X"28",X"14",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"EA",
		X"7A",X"55",X"55",X"95",X"2A",X"54",X"95",X"AA",X"56",X"A1",X"2A",X"55",X"A9",X"5A",X"55",X"AD",
		X"AA",X"54",X"55",X"55",X"55",X"55",X"55",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"55",X"55",
		X"55",X"55",X"55",X"A9",X"AA",X"55",X"AF",X"2A",X"55",X"A9",X"5A",X"55",X"AA",X"56",X"D5",X"AA",
		X"54",X"95",X"AA",X"AA",X"AA",X"AA",X"2A",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"5A",X"95",X"AA",X"AA",X"6A",X"55",X"A5",X"2A",X"55",X"A9",X"5A",X"D5",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"94",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"D4",X"AA",X"AA",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AA",X"56",X"AD",X"6A",X"95",X"AA",X"54",
		X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"C2",X"71",X"87",X"63",X"1C",X"8E",X"E3",X"19",X"8F",X"33",X"E1",X"31",X"1E",X"E3",
		X"71",X"8C",X"E3",X"45",X"E7",X"32",X"57",X"55",X"AA",X"B8",X"8E",X"59",X"E3",X"51",X"55",X"E3",
		X"B8",X"98",X"19",X"57",X"54",X"8D",X"A3",X"2A",X"55",X"2B",X"47",X"AD",X"1A",X"F3",X"18",X"C7",
		X"A3",X"16",X"C7",X"33",X"96",X"E3",X"8C",X"AB",X"C6",X"45",X"57",X"95",X"3C",X"AE",X"B3",X"CC",
		X"71",X"1C",X"C7",X"71",X"9A",X"8B",X"D3",X"E4",X"58",X"B5",X"E2",X"70",X"9C",X"71",X"1C",X"C7",
		X"31",X"4A",X"95",X"0E",X"47",X"A5",X"1A",X"A7",X"2A",X"47",X"93",X"AA",X"B2",X"4C",X"0D",X"C7",
		X"E1",X"AA",X"2A",X"15",X"47",X"2D",X"8E",X"A3",X"70",X"1C",X"E3",X"70",X"38",X"1E",X"57",X"AA",
		X"D6",X"B9",X"5A",X"9D",X"C7",X"D5",X"E9",X"75",X"F5",X"F5",X"FA",X"EC",X"7A",X"5E",X"5D",X"3D",
		X"8E",X"8E",X"A6",X"5C",X"1C",X"97",X"AA",X"AB",X"5A",X"15",X"84",X"81",X"50",X"94",X"42",X"E1",
		X"60",X"70",X"3A",X"5D",X"8B",X"02",X"10",X"0A",X"57",X"4B",X"11",X"89",X"53",X"BF",X"CF",X"87",
		X"01",X"8C",X"D6",X"57",X"97",X"A2",X"A2",X"57",X"FF",X"F5",X"62",X"60",X"78",X"7C",X"9E",X"AE",
		X"70",X"F0",X"F8",X"7E",X"BD",X"C2",X"40",X"D1",X"E7",X"D3",X"A1",X"30",X"BD",X"BA",X"DD",X"B7",
		X"30",X"90",X"AA",X"D7",X"D3",X"90",X"A2",X"CB",X"EB",X"D5",X"77",X"61",X"A0",X"78",X"77",X"15",
		X"21",X"AA",X"D5",X"C7",X"D3",X"F3",X"C1",X"C1",X"E1",X"73",X"15",X"0A",X"56",X"E9",X"78",X"F1",
		X"FA",X"02",X"03",X"87",X"4F",X"1D",X"58",X"F0",X"A8",X"2B",X"1B",X"5F",X"1F",X"0C",X"38",X"76",
		X"AB",X"42",X"C1",X"4B",X"D3",X"E1",X"F5",X"7D",X"60",X"E0",X"F0",X"AB",X"0A",X"54",X"BD",X"B8",
		X"62",X"D7",X"F7",X"80",X"81",X"C7",X"1F",X"15",X"8A",X"5E",X"F1",X"E2",X"D5",X"FB",X"02",X"05",
		X"9E",X"7E",X"91",X"A0",X"55",X"3F",X"78",X"F0",X"EB",X"0F",X"38",X"F0",X"F1",X"83",X"0A",X"76",
		X"8B",X"17",X"AE",X"EE",X"3E",X"60",X"C0",X"E7",X"07",X"15",X"F2",X"C5",X"8B",X"CA",X"BB",X"7B",
		X"C0",X"81",X"8F",X"2F",X"48",X"D1",X"57",X"B1",X"C3",X"57",X"7F",X"80",X"81",X"1F",X"3F",X"20",
		X"A5",X"2F",X"DC",X"E0",X"57",X"7F",X"C0",X"80",X"9F",X"57",X"A0",X"D4",X"17",X"AE",X"E8",X"5B",
		X"1F",X"E0",X"C0",X"8F",X"57",X"C0",X"AA",X"17",X"7A",X"D8",X"A7",X"1F",X"70",X"E0",X"17",X"4F",
		X"A0",X"53",X"0F",X"3E",X"F1",X"AB",X"0B",X"38",X"F8",X"C5",X"05",X"E8",X"AA",X"8B",X"47",X"3F",
		X"F5",X"80",X"03",X"7F",X"B4",X"02",X"5E",X"F9",X"E0",X"C5",X"8F",X"0F",X"70",X"F0",X"97",X"AA",
		X"40",X"8F",X"1E",X"76",X"FA",X"F2",X"00",X"07",X"7F",X"AA",X"0A",X"EC",X"D4",X"45",X"97",X"9F",
		X"1E",X"E0",X"E0",X"AF",X"48",X"85",X"2E",X"55",X"BE",X"F4",X"A3",X"01",X"1E",X"7D",X"1A",X"49",
		X"B1",X"A3",X"53",X"57",X"5F",X"0B",X"E0",X"E2",X"57",X"45",X"85",X"AE",X"E8",X"55",X"5F",X"AD",
		X"00",X"D5",X"8B",X"5D",X"A8",X"54",X"A9",X"5E",X"F5",X"6A",X"03",X"55",X"AA",X"A3",X"55",X"54",
		X"A3",X"AA",X"56",X"D5",X"E9",X"0A",X"55",X"55",X"AA",X"4A",X"55",X"C5",X"AA",X"6A",X"95",X"2A",
		X"D5",X"AA",X"57",X"AC",X"42",X"A5",X"4A",X"B5",X"AA",X"55",X"91",X"AA",X"AA",X"0F",X"55",X"75",
		X"A2",X"AA",X"6A",X"51",X"55",X"54",X"AB",X"AA",X"46",X"55",X"B5",X"AA",X"52",X"A5",X"6A",X"A5",
		X"AA",X"55",X"AA",X"54",X"B5",X"5A",X"95",X"AA",X"55",X"55",X"AA",X"AA",X"78",X"55",X"15",X"AD",
		X"AA",X"2A",X"55",X"55",X"A9",X"AA",X"4A",X"55",X"AD",X"2A",X"55",X"BA",X"56",X"A9",X"5A",X"A5",
		X"6A",X"95",X"AA",X"55",X"A5",X"6A",X"57",X"55",X"55",X"95",X"AA",X"AA",X"54",X"55",X"95",X"B3",
		X"AA",X"4B",X"55",X"55",X"AD",X"AA",X"12",X"D5",X"AA",X"55",X"A9",X"5A",X"95",X"5A",X"55",X"AB",
		X"52",X"95",X"AA",X"6A",X"55",X"55",X"55",X"A4",X"AA",X"2E",X"55",X"55",X"D5",X"AA",X"AA",X"5C",
		X"55",X"A5",X"6A",X"55",X"AA",X"55",X"55",X"55",X"55",X"55",X"55",X"A9",X"8A",X"55",X"55",X"95",
		X"AA",X"AA",X"AA",X"52",X"55",X"55",X"B5",X"AA",X"2A",X"56",X"55",X"AD",X"AA",X"42",X"55",X"AB",
		X"54",X"A7",X"5A",X"55",X"2A",X"55",X"AD",X"4A",X"55",X"8D",X"AA",X"AA",X"55",X"55",X"D6",X"8A",
		X"AA",X"53",X"55",X"95",X"2B",X"AA",X"4E",X"55",X"D5",X"A1",X"2A",X"55",X"EA",X"54",X"AD",X"4A",
		X"95",X"EA",X"55",X"A9",X"55",X"AC",X"78",X"51",X"AB",X"AA",X"0E",X"55",X"55",X"B5",X"A2",X"E8",
		X"53",X"55",X"55",X"D5",X"8B",X"AA",X"AA",X"54",X"55",X"75",X"AD",X"EE",X"56",X"01",X"A8",X"57",
		X"A8",X"5A",X"B5",X"FF",X"55",X"00",X"F0",X"3B",X"4A",X"27",X"22",X"F5",X"BB",X"BB",X"11",X"80",
		X"FD",X"AA",X"AA",X"08",X"6A",X"DF",X"BD",X"2B",X"00",X"F8",X"57",X"55",X"29",X"50",X"BD",X"BB",
		X"DD",X"05",X"00",X"FF",X"2A",X"B5",X"08",X"72",X"EB",X"DB",X"5D",X"01",X"E0",X"EF",X"52",X"15",
		X"41",X"ED",X"AE",X"BB",X"1B",X"00",X"F4",X"AF",X"AA",X"42",X"D0",X"6E",X"F5",X"BE",X"06",X"80",
		X"EE",X"B5",X"AA",X"40",X"B4",X"5B",X"BD",X"AF",X"03",X"40",X"F7",X"55",X"95",X"02",X"FA",X"56",
		X"DD",X"6F",X"01",X"A0",X"5F",X"A7",X"2A",X"90",X"BA",X"5B",X"ED",X"D7",X"00",X"D0",X"AF",X"AB",
		X"4A",X"40",X"B7",X"A9",X"7F",X"57",X"00",X"B0",X"DF",X"55",X"0A",X"44",X"BB",X"D6",X"BD",X"AB",
		X"00",X"D0",X"BF",X"2A",X"45",X"44",X"BB",X"5B",X"DD",X"BB",X"00",X"D0",X"BF",X"52",X"25",X"48",
		X"F7",X"AA",X"DE",X"5D",X"00",X"E8",X"AF",X"AA",X"12",X"44",X"DF",X"A5",X"EE",X"3B",X"00",X"D8",
		X"B7",X"AA",X"0A",X"52",X"ED",X"6A",X"FD",X"AE",X"00",X"B0",X"5F",X"55",X"2A",X"44",X"ED",X"6B",
		X"DD",X"2F",X"00",X"E8",X"6F",X"29",X"15",X"44",X"F7",X"AA",X"FE",X"2E",X"00",X"B8",X"6F",X"55",
		X"25",X"40",X"EF",X"5A",X"FD",X"AE",X"00",X"D0",X"DF",X"52",X"15",X"44",X"BB",X"EA",X"FA",X"5D",
		X"00",X"E0",X"EF",X"52",X"55",X"84",X"EA",X"76",X"ED",X"7B",X"00",X"A0",X"7F",X"95",X"2A",X"41",
		X"EA",X"57",X"DD",X"BB",X"00",X"C0",X"7F",X"55",X"54",X"11",X"EA",X"7A",X"EB",X"7D",X"01",X"80",
		X"FF",X"4A",X"A9",X"12",X"D4",X"FA",X"75",X"BB",X"02",X"00",X"FF",X"AB",X"A8",X"14",X"51",X"ED",
		X"BB",X"DB",X"05",X"00",X"FC",X"AF",X"54",X"2A",X"42",X"B5",X"7F",X"DD",X"05",X"00",X"EC",X"DF",
		X"52",X"15",X"21",X"AA",X"FF",X"5D",X"55",X"00",X"E0",X"DF",X"95",X"4A",X"11",X"A2",X"F7",X"EF",
		X"2A",X"01",X"40",X"EF",X"57",X"55",X"91",X"88",X"DA",X"FF",X"5D",X"04",X"80",X"EA",X"77",X"55",
		X"15",X"22",X"D2",X"FD",X"BF",X"12",X"00",X"A4",X"77",X"B7",X"AA",X"10",X"91",X"FA",X"7F",X"97",
		X"00",X"A0",X"BA",X"DD",X"D5",X"12",X"22",X"6A",X"FD",X"BF",X"0A",X"40",X"A4",X"7A",X"77",X"AB",
		X"44",X"84",X"EA",X"FF",X"AD",X"08",X"20",X"AA",X"DB",X"5D",X"55",X"84",X"A8",X"FA",X"7F",X"55",
		X"04",X"A0",X"6A",X"7D",X"AB",X"55",X"88",X"48",X"FD",X"EF",X"4A",X"10",X"88",X"BA",X"76",X"5D",
		X"95",X"88",X"A8",X"DD",X"7F",X"95",X"20",X"48",X"D5",X"BA",X"75",X"A5",X"48",X"A5",X"DA",X"DF",
		X"AB",X"82",X"20",X"52",X"5D",X"75",X"6D",X"A5",X"88",X"A8",X"FD",X"77",X"55",X"20",X"88",X"4A",
		X"BD",X"BE",X"55",X"0A",X"14",X"AD",X"FF",X"5D",X"25",X"00",X"52",X"75",X"AF",X"AB",X"4A",X"44",
		X"B2",X"FA",X"7F",X"55",X"01",X"20",X"AA",X"D7",X"AB",X"4B",X"45",X"22",X"D5",X"FB",X"5E",X"57",
		X"01",X"20",X"6A",X"77",X"57",X"AB",X"22",X"42",X"D5",X"FB",X"76",X"5D",X"09",X"00",X"D4",X"FB",
		X"56",X"95",X"4A",X"41",X"AA",X"DF",X"AB",X"EA",X"AE",X"00",X"50",X"FD",X"55",X"A9",X"BA",X"08",
		X"51",X"F7",X"B5",X"AA",X"EE",X"0B",X"00",X"55",X"AF",X"55",X"B5",X"5A",X"80",X"EA",X"5D",X"AB",
		X"5A",X"DF",X"8A",X"00",X"69",X"55",X"AB",X"BA",X"0A",X"11",X"F5",X"AA",X"AA",X"5D",X"F7",X"2D",
		X"00",X"A8",X"75",X"AB",X"55",X"2B",X"10",X"B5",X"6F",X"95",X"EA",X"DB",X"5D",X"04",X"40",X"EB",
		X"BA",X"AA",X"54",X"44",X"D5",X"B7",X"8A",X"AA",X"6F",X"DF",X"11",X"00",X"EA",X"5D",X"AB",X"4A",
		X"81",X"AA",X"BD",X"2A",X"56",X"B7",X"FE",X"15",X"00",X"F8",X"AE",X"AA",X"55",X"04",X"D5",X"BE",
		X"4A",X"55",X"D5",X"FE",X"3B",X"00",X"D0",X"EB",X"52",X"97",X"08",X"D5",X"7A",X"55",X"AA",X"54",
		X"FD",X"BF",X"02",X"00",X"77",X"5D",X"AD",X"88",X"A8",X"6E",X"55",X"45",X"55",X"FD",X"FE",X"0B",
		X"00",X"F4",X"EE",X"5A",X"28",X"48",X"DD",X"2E",X"95",X"AA",X"D4",X"FF",X"AE",X"00",X"C0",X"7D",
		X"57",X"85",X"88",X"EA",X"AE",X"52",X"51",X"D5",X"BE",X"BF",X"02",X"00",X"FD",X"5B",X"95",X"08",
		X"D2",X"BB",X"15",X"D1",X"4A",X"F5",X"BF",X"2B",X"00",X"70",X"7F",X"55",X"22",X"A2",X"EE",X"55",
		X"11",X"55",X"AD",X"FE",X"5B",X"05",X"00",X"EF",X"57",X"89",X"50",X"B5",X"6E",X"15",X"8A",X"56",
		X"EF",X"FE",X"4A",X"00",X"F0",X"6F",X"A9",X"08",X"6A",X"5F",X"55",X"14",X"A9",X"BB",X"BB",X"57",
		X"05",X"80",X"BF",X"55",X"23",X"50",X"ED",X"55",X"A9",X"48",X"F5",X"AB",X"FD",X"55",X"00",X"F8",
		X"BA",X"AA",X"40",X"F4",X"55",X"D1",X"8A",X"E8",X"5E",X"DD",X"BD",X"00",X"60",X"DF",X"AA",X"05",
		X"A8",X"77",X"A5",X"4A",X"A4",X"BB",X"D5",X"DF",X"12",X"80",X"F8",X"5B",X"55",X"40",X"ED",X"AA",
		X"8B",X"A0",X"7D",X"55",X"FF",X"8A",X"02",X"44",X"BF",X"4B",X"11",X"AA",X"5D",X"AA",X"14",X"B8",
		X"57",X"F5",X"AF",X"A8",X"00",X"DC",X"57",X"A5",X"A0",X"EA",X"56",X"15",X"50",X"5F",X"A9",X"7F",
		X"55",X"01",X"D0",X"3F",X"55",X"0A",X"72",X"BB",X"52",X"85",X"EA",X"55",X"FB",X"AB",X"1A",X"00",
		X"FD",X"95",X"2A",X"42",X"DB",X"15",X"17",X"D0",X"BB",X"AA",X"5F",X"55",X"01",X"68",X"5F",X"39",
		X"12",X"EC",X"56",X"B5",X"48",X"D5",X"AA",X"F7",X"5D",X"15",X"80",X"FA",X"AA",X"45",X"50",X"57",
		X"55",X"2B",X"A8",X"7A",X"75",X"77",X"57",X"01",X"A8",X"5F",X"B5",X"00",X"F5",X"AA",X"54",X"A1",
		X"5A",X"A7",X"7E",X"57",X"1D",X"80",X"BA",X"AB",X"03",X"54",X"57",X"D5",X"0A",X"F8",X"4A",X"F5",
		X"EB",X"AA",X"01",X"74",X"AB",X"5E",X"80",X"76",X"A5",X"2B",X"01",X"BF",X"54",X"BF",X"AA",X"2B",
		X"80",X"57",X"D5",X"07",X"D8",X"2A",X"FA",X"02",X"75",X"45",X"F7",X"D6",X"AE",X"02",X"B8",X"74",
		X"BB",X"40",X"B5",X"D2",X"15",X"AA",X"56",X"EA",X"5B",X"5F",X"15",X"C0",X"AA",X"EB",X"0A",X"54",
		X"55",X"7D",X"09",X"B8",X"8B",X"7E",X"5B",X"57",X"01",X"AA",X"7A",X"17",X"60",X"55",X"AD",X"55",
		X"A0",X"AE",X"F4",X"BA",X"5B",X"0D",X"C0",X"A5",X"AF",X"0A",X"AA",X"52",X"77",X"11",X"F4",X"89",
		X"AF",X"BB",X"BA",X"00",X"56",X"ED",X"56",X"A0",X"AA",X"DC",X"89",X"42",X"8F",X"3E",X"FD",X"AA",
		X"03",X"B0",X"74",X"57",X"21",X"2E",X"5A",X"57",X"54",X"E8",X"A3",X"77",X"57",X"17",X"C0",X"52",
		X"BF",X"02",X"55",X"AA",X"57",X"B4",X"42",X"97",X"EE",X"BE",X"55",X"01",X"2C",X"FD",X"2A",X"A8",
		X"A2",X"5D",X"55",X"15",X"B5",X"EC",X"EB",X"6B",X"05",X"50",X"F4",X"AB",X"14",X"29",X"56",X"2F",
		X"4A",X"55",X"EA",X"DD",X"B7",X"0A",X"A0",X"F0",X"57",X"15",X"89",X"AA",X"76",X"05",X"9D",X"E8",
		X"DE",X"7D",X"55",X"80",X"C2",X"5F",X"95",X"42",X"55",X"BA",X"07",X"AE",X"70",X"DD",X"FA",X"AA",
		X"01",X"06",X"F7",X"55",X"89",X"2A",X"BA",X"5A",X"F0",X"41",X"1F",X"EF",X"AA",X"03",X"0C",X"FC",
		X"AA",X"15",X"B4",X"70",X"97",X"2A",X"5C",X"E9",X"76",X"77",X"09",X"28",X"F8",X"EA",X"15",X"51",
		X"D1",X"D5",X"16",X"BA",X"E0",X"D3",X"5F",X"5D",X"A0",X"A0",X"CB",X"37",X"68",X"C1",X"AA",X"D5",
		X"C1",X"43",X"D7",X"EE",X"EA",X"01",X"03",X"8F",X"AF",X"E2",X"82",X"43",X"4F",X"55",X"A5",X"AA",
		X"EB",X"6B",X"0B",X"04",X"4D",X"BB",X"4B",X"07",X"86",X"47",X"8F",X"47",X"A3",X"EB",X"D5",X"07",
		X"0E",X"38",X"7A",X"D5",X"05",X"07",X"97",X"8D",X"AB",X"AA",X"F2",X"D5",X"73",X"50",X"70",X"E8",
		X"7A",X"39",X"12",X"95",X"2E",X"F2",X"E8",X"72",X"BD",X"AE",X"A8",X"40",X"D1",X"D5",X"A7",X"8A",
		X"8A",X"5A",X"55",X"97",X"AA",X"7A",X"7D",X"1D",X"06",X"0C",X"76",X"BD",X"38",X"54",X"2A",X"55",
		X"C7",X"C3",X"E5",X"EA",X"7A",X"70",X"50",X"98",X"D5",X"E3",X"A1",X"A1",X"CA",X"72",X"79",X"59",
		X"5D",X"B7",X"8B",X"82",X"82",X"55",X"AF",X"0E",X"95",X"8A",X"16",X"2F",X"1E",X"DD",X"EA",X"6B",
		X"70",X"50",X"34",X"3E",X"7A",X"38",X"54",X"CC",X"AC",X"BA",X"CA",X"D5",X"75",X"87",X"83",X"C2",
		X"D1",X"A3",X"47",X"83",X"C3",X"C5",X"AA",X"5D",X"AD",X"AE",X"2B",X"1C",X"14",X"56",X"5D",X"3D",
		X"3C",X"38",X"38",X"7A",X"78",X"3C",X"3E",X"5D",X"71",X"30",X"38",X"56",X"ED",X"E2",X"50",X"A9",
		X"38",X"9D",X"AE",X"56",X"D7",X"8B",X"02",X"15",X"1D",X"8F",X"8F",X"26",X"15",X"55",X"3E",X"AE",
		X"5A",X"57",X"7D",X"38",X"18",X"38",X"75",X"7A",X"74",X"A8",X"68",X"9C",X"4E",X"57",X"D7",X"E9",
		X"E1",X"C0",X"E0",X"D4",X"D5",X"C5",X"A2",X"A2",X"AA",X"3A",X"5D",X"57",X"57",X"07",X"07",X"83",
		X"AA",X"1E",X"8F",X"0E",X"45",X"8B",X"97",X"C7",X"E3",X"D5",X"2B",X"0C",X"06",X"57",X"AD",X"AE",
		X"8A",X"52",X"55",X"BC",X"AA",X"AE",X"5D",X"5D",X"31",X"28",X"18",X"B7",X"EA",X"54",X"A4",X"54",
		X"D5",X"EA",X"D5",X"BA",X"EE",X"E1",X"40",X"70",X"74",X"D5",X"A3",X"A2",X"E2",X"F0",X"71",X"55",
		X"5D",X"B7",X"83",X"83",X"C2",X"D1",X"B3",X"C3",X"91",X"AA",X"54",X"3D",X"4E",X"DD",X"BA",X"0E",
		X"07",X"86",X"A6",X"AB",X"4E",X"14",X"95",X"A9",X"B3",X"71",X"71",X"F7",X"6A",X"38",X"50",X"B4",
		X"BA",X"55",X"2A",X"52",X"85",X"C7",X"C7",X"E3",X"5A",X"5F",X"31",X"A0",X"A8",X"AE",X"AB",X"11",
		X"15",X"1D",X"1F",X"2E",X"8E",X"77",X"F5",X"44",X"01",X"87",X"8F",X"17",X"87",X"52",X"A5",X"E3",
		X"65",X"A9",X"DC",X"9D",X"0F",X"0C",X"34",X"76",X"AB",X"2A",X"52",X"74",X"55",X"1E",X"3A",X"5E",
		X"5D",X"5F",X"A0",X"A0",X"D2",X"AF",X"4A",X"85",X"AA",X"55",X"C3",X"C3",X"E3",X"EB",X"7C",X"0A",
		X"01",X"C7",X"DD",X"AA",X"A8",X"B0",X"56",X"1D",X"1E",X"36",X"ED",X"EB",X"A3",X"20",X"F0",X"F4",
		X"AA",X"54",X"A4",X"5A",X"75",X"E2",X"70",X"B9",X"7B",X"3D",X"81",X"82",X"47",X"5F",X"51",X"51",
		X"A9",X"6B",X"0A",X"17",X"57",X"EF",X"E3",X"03",X"14",X"7C",X"EA",X"45",X"25",X"16",X"BD",X"2A",
		X"95",X"AA",X"5E",X"5F",X"AB",X"80",X"81",X"D7",X"5B",X"D0",X"D0",X"A5",X"1B",X"AA",X"A2",X"A7",
		X"6F",X"75",X"05",X"14",X"BA",X"EB",X"42",X"15",X"B9",X"DA",X"05",X"2B",X"D5",X"E5",X"4F",X"5F",
		X"40",X"81",X"1F",X"7D",X"50",X"43",X"8F",X"AE",X"50",X"87",X"AF",X"7A",X"D5",X"2A",X"70",X"F0",
		X"A9",X"0D",X"6A",X"D4",X"A5",X"2E",X"78",X"D1",X"4D",X"BF",X"EC",X"02",X"03",X"5F",X"D5",X"05",
		X"4D",X"BA",X"A6",X"2A",X"7C",X"F0",X"55",X"1F",X"BD",X"C0",X"41",X"9F",X"5C",X"C1",X"43",X"57",
		X"A9",X"51",X"4D",X"FA",X"F4",X"C5",X"07",X"B8",X"E0",X"47",X"17",X"D4",X"54",X"5D",X"B4",X"A2",
		X"8B",X"BE",X"7A",X"55",X"05",X"16",X"FA",X"54",X"07",X"2E",X"D5",X"A9",X"5A",X"E8",X"E2",X"5D",
		X"AF",X"6A",X"C0",X"81",X"1F",X"DD",X"A0",X"26",X"3D",X"55",X"15",X"AE",X"EC",X"D6",X"55",X"17",
		X"B0",X"F0",X"C5",X"2E",X"70",X"A1",X"57",X"B1",X"C2",X"87",X"BE",X"BA",X"55",X"03",X"16",X"BE",
		X"AA",X"0A",X"3A",X"F4",X"45",X"1D",X"5C",X"E9",X"AE",X"AE",X"5A",X"40",X"45",X"9F",X"6A",X"41",
		X"2B",X"5E",X"D1",X"0A",X"57",X"EA",X"6B",X"D7",X"0A",X"A8",X"D8",X"57",X"15",X"B4",X"A2",X"17",
		X"55",X"D1",X"A5",X"BE",X"6E",X"55",X"01",X"2B",X"7A",X"D5",X"82",X"56",X"EC",X"62",X"15",X"BA",
		X"D4",X"AF",X"AE",X"3A",X"C0",X"C1",X"57",X"35",X"A2",X"8E",X"BA",X"A8",X"45",X"5D",X"7C",X"ED",
		X"AA",X"0A",X"2C",X"F4",X"D1",X"0B",X"74",X"E2",X"53",X"95",X"AA",X"55",X"AF",X"5E",X"55",X"A0",
		X"8A",X"9E",X"76",X"44",X"95",X"BA",X"A2",X"13",X"5D",X"BC",X"AB",X"AB",X"07",X"54",X"A8",X"4F",
		X"55",X"AA",X"54",X"AB",X"54",X"A5",X"AA",X"DD",X"AD",X"BE",X"00",X"0B",X"7E",X"D4",X"05",X"9D",
		X"F8",X"C2",X"86",X"5E",X"F4",X"55",X"5D",X"15",X"A8",X"AA",X"53",X"55",X"D1",X"4A",X"17",X"3A",
		X"5A",X"B5",X"6E",X"B5",X"AB",X"40",X"89",X"5E",X"55",X"29",X"56",X"7C",X"A8",X"45",X"5D",X"75",
		X"57",X"BB",X"0A",X"58",X"D4",X"55",X"55",X"D4",X"8A",X"AA",X"AA",X"AA",X"5D",X"7D",X"75",X"03",
		X"B8",X"F0",X"45",X"17",X"6A",X"55",X"2D",X"5A",X"B1",X"AA",X"57",X"AB",X"5B",X"90",X"2A",X"55",
		X"A9",X"4A",X"D5",X"AA",X"54",X"55",X"D5",X"AA",X"AF",X"2E",X"14",X"54",X"55",X"87",X"96",X"AA",
		X"AA",X"2A",X"5A",X"55",X"DD",X"97",X"BE",X"E0",X"A0",X"13",X"5D",X"B1",X"8A",X"55",X"AA",X"55",
		X"A5",X"5A",X"BD",X"EA",X"45",X"07",X"2E",X"74",X"A9",X"54",X"E9",X"8A",X"56",X"55",X"55",X"BD",
		X"AA",X"2F",X"3C",X"70",X"51",X"47",X"AE",X"A8",X"2A",X"1B",X"75",X"D1",X"45",X"9F",X"EA",X"8A",
		X"17",X"AC",X"52",X"95",X"AA",X"54",X"A5",X"1A",X"5D",X"EA",X"54",X"AF",X"5A",X"55",X"05",X"AB",
		X"E8",X"A2",X"16",X"5D",X"54",X"15",X"2F",X"EA",X"E2",X"8B",X"5E",X"D1",X"45",X"95",X"AA",X"AA",
		X"4A",X"55",X"AA",X"54",X"B5",X"4A",X"9D",X"EA",X"55",X"AB",X"5A",X"51",X"2A",X"55",X"A9",X"62",
		X"55",X"AB",X"AA",X"54",X"55",X"57",X"D5",X"AA",X"AA",X"A8",X"54",X"55",X"55",X"51",X"AB",X"AA",
		X"AA",X"6A",X"55",X"55",X"AD",X"AA",X"2A",X"55",X"AA",X"56",X"A9",X"52",X"D5",X"2A",X"55",X"55",
		X"55",X"D5",X"AA",X"56",X"55",X"A9",X"AA",X"AA",X"60",X"55",X"55",X"55",X"A9",X"AA",X"AA",X"FA",
		X"54",X"55",X"55",X"55",X"AA",X"AA",X"2A",X"55",X"AD",X"4A",X"D5",X"AA",X"54",X"AD",X"52",X"95",
		X"AA",X"55",X"AB",X"52",X"95",X"AA",X"56",X"55",X"55",X"AB",X"AA",X"AA",X"55",X"A9",X"AA",X"AA",
		X"B5",X"29",X"55",X"BD",X"5B",X"AB",X"10",X"A5",X"A4",X"2A",X"25",X"A9",X"AA",X"AA",X"6A",X"DF",
		X"6E",X"AD",X"AA",X"54",X"25",X"A2",X"22",X"49",X"4A",X"A9",X"AA",X"DB",X"DB",X"AA",X"12",X"A5",
		X"AA",X"BA",X"6E",X"BB",X"AA",X"A2",X"52",X"25",X"A2",X"4A",X"55",X"B5",X"DA",X"A5",X"AE",X"AD",
		X"4A",X"55",X"55",X"AA",X"5A",X"DF",X"5D",X"55",X"24",X"29",X"52",X"A5",X"DA",X"6E",X"57",X"A5",
		X"A4",X"88",X"24",X"29",X"B5",X"B6",X"5D",X"A9",X"AA",X"4B",X"52",X"B5",X"F6",X"55",X"A9",X"EA",
		X"AD",X"02",X"92",X"AA",X"AA",X"5A",X"EF",X"EE",X"AA",X"20",X"55",X"4A",X"49",X"55",X"D5",X"DD",
		X"56",X"21",X"A5",X"AA",X"44",X"48",X"52",X"ED",X"5B",X"AD",X"7D",X"DB",X"5A",X"A9",X"A2",X"4A",
		X"A9",X"92",X"48",X"A9",X"76",X"DF",X"AA",X"B6",X"AB",X"22",X"22",X"A9",X"AA",X"48",X"A9",X"6A",
		X"DB",X"57",X"AB",X"0A",X"55",X"AA",X"2A",X"51",X"AA",X"6A",X"AD",X"4A",X"D5",X"FE",X"DB",X"56",
		X"6B",X"AB",X"84",X"10",X"AA",X"4A",X"55",X"55",X"ED",X"DD",X"2A",X"48",X"A5",X"94",X"44",X"52",
		X"F7",X"6D",X"BB",X"D5",X"AA",X"82",X"24",X"91",X"AA",X"AA",X"55",X"95",X"52",X"F7",X"56",X"A4",
		X"F5",X"BB",X"2A",X"91",X"AA",X"A4",X"12",X"55",X"75",X"AF",X"22",X"92",X"D4",X"B6",X"5B",X"BB",
		X"B5",X"4B",X"40",X"20",X"A9",X"B6",X"5B",X"AB",X"DE",X"B7",X"0A",X"82",X"D4",X"5E",X"09",X"A4",
		X"FA",X"56",X"21",X"A9",X"BF",X"AB",X"04",X"A2",X"DA",X"DE",X"2A",X"E9",X"6D",X"9B",X"40",X"54",
		X"BF",X"B5",X"90",X"54",X"AB",X"55",X"08",X"C9",X"FE",X"5F",X"09",X"D2",X"FE",X"4A",X"00",X"D4",
		X"BE",X"15",X"20",X"DD",X"6F",X"09",X"52",X"EF",X"BB",X"00",X"20",X"DB",X"5B",X"21",X"E9",X"FF",
		X"2B",X"20",X"BA",X"7F",X"05",X"A0",X"BA",X"AF",X"02",X"A1",X"F6",X"5B",X"21",X"54",X"F7",X"56",
		X"08",X"D9",X"FF",X"15",X"40",X"EA",X"DF",X"04",X"48",X"FB",X"B7",X"82",X"A8",X"BB",X"25",X"20",
		X"E9",X"FF",X"4E",X"40",X"FA",X"5F",X"01",X"80",X"FE",X"2B",X"00",X"ED",X"FF",X"09",X"A0",X"FE",
		X"2D",X"40",X"DA",X"B7",X"52",X"92",X"F5",X"BD",X"05",X"00",X"EF",X"AF",X"00",X"A4",X"FF",X"17",
		X"00",X"FD",X"5F",X"00",X"D0",X"7F",X"8B",X"20",X"F5",X"DD",X"92",X"40",X"FE",X"DF",X"00",X"C0",
		X"FF",X"0F",X"00",X"FC",X"7F",X"01",X"A8",X"FF",X"15",X"00",X"FC",X"FF",X"00",X"60",X"FF",X"2F",
		X"00",X"E8",X"FF",X"01",X"80",X"FF",X"3F",X"00",X"F8",X"FF",X"01",X"80",X"FF",X"0F",X"00",X"FD",
		X"5F",X"01",X"A0",X"FF",X"4F",X"00",X"F8",X"FF",X"01",X"80",X"FF",X"1F",X"00",X"FC",X"7F",X"00",
		X"F0",X"FF",X"03",X"C0",X"FF",X"0B",X"00",X"ED",X"BF",X"02",X"80",X"FF",X"9F",X"00",X"F0",X"FF",
		X"01",X"C0",X"FF",X"07",X"00",X"FF",X"1F",X"00",X"FC",X"3F",X"00",X"EC",X"FF",X"00",X"E0",X"FF",
		X"03",X"00",X"FF",X"07",X"00",X"FF",X"1F",X"00",X"FE",X"1F",X"00",X"FC",X"7F",X"00",X"F8",X"FF",
		X"00",X"E0",X"FF",X"01",X"E0",X"FF",X"01",X"E0",X"FF",X"00",X"F8",X"3F",X"00",X"FC",X"1F",X"00",
		X"FE",X"27",X"00",X"FF",X"3F",X"00",X"FC",X"1F",X"00",X"FF",X"07",X"C0",X"FF",X"01",X"F0",X"3F",
		X"00",X"FE",X"07",X"40",X"FF",X"3B",X"00",X"FF",X"07",X"C0",X"FF",X"00",X"F8",X"3F",X"00",X"FE",
		X"07",X"80",X"FF",X"01",X"F0",X"3F",X"00",X"FE",X"0F",X"80",X"FF",X"03",X"F0",X"7F",X"00",X"FC",
		X"1F",X"00",X"FE",X"07",X"C0",X"FF",X"01",X"E0",X"7F",X"00",X"FC",X"4F",X"00",X"FF",X"13",X"C0",
		X"7F",X"07",X"E0",X"FF",X"00",X"F8",X"1F",X"00",X"FF",X"03",X"E0",X"7F",X"00",X"FC",X"1F",X"00",
		X"FF",X"07",X"80",X"FF",X"03",X"E0",X"7F",X"00",X"F8",X"1F",X"00",X"FF",X"03",X"E0",X"FF",X"00",
		X"F8",X"3F",X"00",X"FE",X"0F",X"80",X"FF",X"03",X"E0",X"7F",X"00",X"FE",X"0F",X"80",X"FF",X"01",
		X"E0",X"FF",X"00",X"E0",X"7F",X"00",X"F8",X"1F",X"80",X"FF",X"07",X"C0",X"FF",X"00",X"F8",X"1F",
		X"00",X"FE",X"0F",X"80",X"FF",X"03",X"C0",X"FF",X"01",X"E0",X"FF",X"00",X"F0",X"3F",X"00",X"FF",
		X"07",X"C0",X"FF",X"00",X"F0",X"7F",X"00",X"FC",X"1F",X"00",X"FF",X"03",X"E0",X"FF",X"00",X"FC",
		X"3F",X"00",X"FE",X"0F",X"00",X"FF",X"03",X"E0",X"FF",X"00",X"F8",X"7F",X"00",X"FC",X"1F",X"80",
		X"FF",X"03",X"F0",X"7F",X"00",X"FC",X"0B",X"C0",X"7F",X"02",X"E0",X"FF",X"00",X"F8",X"1F",X"00",
		X"FF",X"07",X"A0",X"FF",X"01",X"F0",X"7F",X"00",X"FC",X"0F",X"C0",X"FF",X"00",X"DC",X"3F",X"60",
		X"E1",X"7F",X"00",X"FC",X"0F",X"80",X"FF",X"03",X"E0",X"FF",X"01",X"F0",X"7F",X"00",X"FC",X"0F",
		X"80",X"FF",X"00",X"E0",X"3F",X"00",X"FE",X"1F",X"00",X"FE",X"07",X"C0",X"FF",X"01",X"F0",X"7F",
		X"00",X"FE",X"13",X"80",X"3F",X"0F",X"E0",X"CF",X"03",X"F8",X"3F",X"00",X"FF",X"0F",X"C0",X"FF",
		X"00",X"E1",X"3F",X"20",X"FC",X"07",X"98",X"7F",X"00",X"FF",X"07",X"E0",X"9F",X"9C",X"A2",X"E7",
		X"1D",X"C0",X"1F",X"0F",X"F0",X"DF",X"01",X"FC",X"0F",X"C0",X"FF",X"00",X"FC",X"07",X"C0",X"3F",
		X"A0",X"FC",X"03",X"C0",X"FF",X"30",X"F0",X"1F",X"00",X"FE",X"07",X"C0",X"FF",X"00",X"F8",X"0F",
		X"A8",X"FF",X"08",X"FC",X"07",X"87",X"E3",X"F0",X"0B",X"E0",X"FF",X"00",X"FC",X"1F",X"80",X"FF",
		X"03",X"C0",X"FF",X"00",X"FC",X"1F",X"00",X"FE",X"03",X"E0",X"7F",X"03",X"E0",X"7F",X"00",X"FE",
		X"07",X"E0",X"7F",X"20",X"F4",X"0F",X"0E",X"F0",X"DF",X"00",X"FE",X"0F",X"E0",X"FF",X"00",X"FE",
		X"1F",X"80",X"F7",X"07",X"C0",X"FF",X"03",X"F0",X"7F",X"00",X"FC",X"07",X"F0",X"7F",X"00",X"FC",
		X"3F",X"00",X"FC",X"1F",X"40",X"FF",X"03",X"F8",X"2F",X"E0",X"75",X"F0",X"1F",X"00",X"FF",X"03",
		X"F8",X"1F",X"80",X"FF",X"01",X"F0",X"3F",X"20",X"7E",X"1C",X"06",X"8F",X"F0",X"79",X"C0",X"7F",
		X"82",X"FE",X"07",X"F8",X"1F",X"C0",X"FF",X"00",X"F8",X"07",X"78",X"7E",X"E0",X"07",X"86",X"3F",
		X"C0",X"FB",X"03",X"F0",X"1F",X"10",X"FC",X"87",X"00",X"FF",X"03",X"E0",X"FF",X"00",X"FE",X"17",
		X"F0",X"8F",X"04",X"FE",X"21",X"C1",X"7F",X"08",X"FC",X"09",X"5D",X"06",X"6F",X"0B",X"E0",X"7F",
		X"00",X"FE",X"03",X"E0",X"FF",X"00",X"FC",X"1F",X"80",X"FF",X"03",X"F8",X"3F",X"00",X"FF",X"07",
		X"E0",X"FF",X"00",X"FE",X"23",X"F0",X"07",X"0D",X"8D",X"CD",X"81",X"F1",X"17",X"52",X"FD",X"B1",
		X"40",X"FF",X"17",X"C0",X"FF",X"01",X"F0",X"3F",X"00",X"FE",X"07",X"E0",X"FF",X"00",X"FC",X"1F",
		X"80",X"FF",X"03",X"F0",X"1F",X"00",X"FF",X"04",X"FA",X"87",X"AB",X"E8",X"FA",X"01",X"F0",X"7F",
		X"00",X"FE",X"07",X"C0",X"BF",X"00",X"FC",X"5B",X"C0",X"3F",X"05",X"FC",X"55",X"C0",X"0F",X"57",
		X"FB",X"80",X"FF",X"01",X"F0",X"1F",X"00",X"FF",X"01",X"F0",X"1F",X"80",X"FF",X"82",X"6A",X"7F",
		X"41",X"DC",X"1F",X"04",X"FF",X"03",X"E2",X"3F",X"60",X"F4",X"05",X"0F",X"7D",X"C1",X"EA",X"0F",
		X"68",X"BF",X"00",X"7F",X"C1",X"F6",X"01",X"F0",X"3F",X"80",X"7F",X"07",X"F8",X"47",X"B9",X"17",
		X"A0",X"3F",X"01",X"F0",X"1F",X"E0",X"FE",X"04",X"EE",X"07",X"C9",X"FF",X"00",X"F5",X"1F",X"00",
		X"FF",X"02",X"C1",X"B7",X"68",X"D0",X"9F",X"04",X"FC",X"17",X"A0",X"FF",X"01",X"FE",X"0F",X"E0",
		X"BF",X"02",X"FC",X"1F",X"80",X"7F",X"02",X"F8",X"8F",X"80",X"FF",X"01",X"EA",X"15",X"2A",X"6D",
		X"5B",X"81",X"FB",X"07",X"F0",X"7F",X"00",X"FE",X"06",X"F0",X"41",X"DD",X"5E",X"C0",X"7F",X"01",
		X"FC",X"0F",X"B0",X"FF",X"00",X"FC",X"0F",X"80",X"FF",X"01",X"FC",X"1F",X"80",X"FF",X"01",X"D8",
		X"BF",X"80",X"EA",X"5F",X"80",X"FE",X"03",X"F0",X"1F",X"11",X"FE",X"40",X"5F",X"13",X"F4",X"45",
		X"A4",X"3F",X"80",X"FD",X"03",X"C0",X"FF",X"02",X"F8",X"FF",X"00",X"FC",X"17",X"40",X"FF",X"21",
		X"B9",X"17",X"B4",X"44",X"E9",X"07",X"A0",X"FF",X"81",X"FA",X"1A",X"54",X"F5",X"16",X"40",X"FF",
		X"03",X"E8",X"7F",X"00",X"FE",X"07",X"A0",X"FF",X"00",X"F8",X"3F",X"00",X"FF",X"03",X"F0",X"2F",
		X"24",X"FD",X"81",X"8A",X"9F",X"76",X"80",X"FD",X"07",X"80",X"FF",X"01",X"FC",X"2F",X"00",X"FF",
		X"0B",X"C0",X"FF",X"03",X"64",X"3F",X"40",X"F2",X"1F",X"10",X"FE",X"07",X"84",X"FF",X"00",X"F9",
		X"1F",X"A0",X"FF",X"01",X"F8",X"1F",X"80",X"FF",X"17",X"50",X"DF",X"05",X"A0",X"7F",X"01",X"FD",
		X"17",X"A0",X"EF",X"00",X"FC",X"1F",X"80",X"FF",X"05",X"64",X"5F",X"94",X"E4",X"A9",X"8F",X"2C",
		X"FA",X"03",X"48",X"7F",X"48",X"F5",X"5D",X"81",X"F4",X"1F",X"00",X"FE",X"07",X"D0",X"FF",X"00",
		X"FC",X"0F",X"80",X"FF",X"01",X"F0",X"3F",X"00",X"FC",X"0F",X"80",X"FF",X"03",X"F0",X"7F",X"01",
		X"B9",X"7F",X"00",X"FA",X"0F",X"80",X"FF",X"01",X"F0",X"3F",X"00",X"FF",X"03",X"F0",X"7F",X"01",
		X"FA",X"2F",X"40",X"B6",X"1F",X"81",X"F6",X"8F",X"80",X"FE",X"2B",X"C0",X"BF",X"02",X"FC",X"4B",
		X"A0",X"5F",X"29",X"70",X"B7",X"05",X"B8",X"B7",X"00",X"FD",X"2B",X"A8",X"FD",X"81",X"2A",X"3F",
		X"A8",X"ED",X"07",X"AA",X"5F",X"01",X"F7",X"02",X"F4",X"3E",X"90",X"55",X"0F",X"F2",X"93",X"A2",
		X"FC",X"00",X"DB",X"1F",X"F0",X"5B",X"01",X"FF",X"07",X"F0",X"5F",X"01",X"FC",X"0F",X"E0",X"5F",
		X"0A",X"78",X"97",X"02",X"BF",X"15",X"C0",X"5F",X"05",X"F8",X"3F",X"00",X"FF",X"07",X"E0",X"5F",
		X"40",X"FA",X"0B",X"49",X"FF",X"20",X"ED",X"5E",X"A4",X"2A",X"E5",X"05",X"54",X"FB",X"02",X"DA",
		X"1F",X"D0",X"FF",X"00",X"FA",X"1F",X"20",X"ED",X"17",X"40",X"FF",X"01",X"E0",X"FF",X"00",X"F8",
		X"3F",X"00",X"FF",X"07",X"E0",X"7F",X"00",X"F6",X"4B",X"40",X"FD",X"25",X"A0",X"FD",X"0B",X"E0",
		X"FF",X"02",X"F4",X"5F",X"00",X"FB",X"0F",X"80",X"FF",X"02",X"F0",X"3F",X"80",X"FE",X"23",X"A4",
		X"DD",X"4A",X"20",X"EF",X"15",X"C0",X"DF",X"02",X"F4",X"7F",X"00",X"FB",X"1F",X"80",X"FF",X"03",
		X"F0",X"7F",X"00",X"EC",X"1F",X"00",X"FD",X"2B",X"00",X"FF",X"23",X"C0",X"FF",X"09",X"F0",X"BF",
		X"00",X"FE",X"17",X"80",X"FF",X"03",X"E0",X"7F",X"01",X"FC",X"2F",X"80",X"FA",X"17",X"40",X"FF",
		X"05",X"E0",X"7F",X"01",X"FC",X"2F",X"40",X"FF",X"06",X"A0",X"FF",X"03",X"F0",X"7F",X"00",X"FE",
		X"0B",X"A0",X"BF",X"44",X"EA",X"96",X"24",X"DE",X"95",X"A0",X"7F",X"21",X"F4",X"0F",X"A4",X"DE",
		X"0A",X"69",X"DF",X"00",X"EC",X"1E",X"50",X"BB",X"15",X"BA",X"6D",X"A5",X"5A",X"AB",X"AA",X"B4",
		X"52",X"9D",X"12",X"BA",X"17",X"C8",X"B7",X"02",X"FA",X"36",X"48",X"6F",X"2B",X"52",X"FD",X"57",
		X"44",X"7D",X"05",X"F0",X"5B",X"40",X"FF",X"02",X"E8",X"BF",X"00",X"FC",X"2F",X"A0",X"FD",X"03",
		X"E8",X"AF",X"80",X"BA",X"0B",X"A0",X"FB",X"8A",X"F4",X"BB",X"22",X"69",X"B7",X"20",X"EA",X"AF",
		X"80",X"FE",X"07",X"A8",X"BE",X"02",X"EA",X"BB",X"20",X"FA",X"57",X"C8",X"EE",X"12",X"54",X"BD",
		X"02",X"D8",X"5F",X"80",X"FA",X"2B",X"E0",X"DF",X"4A",X"EA",X"D6",X"04",X"D2",X"9D",X"80",X"FE",
		X"15",X"A2",X"5F",X"85",X"F4",X"2D",X"91",X"DA",X"2B",X"48",X"7B",X"91",X"AA",X"AF",X"A0",X"AA",
		X"57",X"2A",X"FD",X"25",X"C1",X"BE",X"10",X"E8",X"2E",X"41",X"F5",X"56",X"E0",X"FF",X"21",X"D8",
		X"57",X"20",X"F7",X"01",X"F0",X"3F",X"81",X"FE",X"07",X"C8",X"BF",X"04",X"EA",X"85",X"B6",X"BA",
		X"B8",X"27",X"5A",X"37",X"C0",X"AD",X"08",X"7C",X"27",X"A4",X"BB",X"44",X"7B",X"4B",X"64",X"55",
		X"A1",X"FD",X"12",X"FD",X"95",X"EA",X"2A",X"00",X"7A",X"81",X"7E",X"83",X"BE",X"7E",X"01",X"FF",
		X"01",X"E0",X"97",X"D0",X"5F",X"41",X"FF",X"82",X"FE",X"01",X"D1",X"2F",X"C0",X"3F",X"01",X"FE",
		X"07",X"E8",X"17",X"A0",X"5B",X"55",X"95",X"52",X"91",X"56",X"FF",X"17",X"B5",X"8B",X"DA",X"50",
		X"45",X"50",X"AF",X"A8",X"D6",X"AD",X"C0",X"BF",X"88",X"24",X"91",X"BC",X"25",X"F4",X"3F",X"FA",
		X"9F",X"00",X"FE",X"02",X"EC",X"03",X"AA",X"7B",X"82",X"FF",X"01",X"B6",X"00",X"F7",X"05",X"E9",
		X"57",X"E0",X"FF",X"02",X"F5",X"0F",X"D0",X"7F",X"22",X"52",X"92",X"56",X"C8",X"FE",X"02",X"59",
		X"2B",X"21",X"6D",X"5F",X"85",X"FE",X"87",X"F0",X"FF",X"00",X"F4",X"03",X"F8",X"07",X"ED",X"6E",
		X"A0",X"77",X"A1",X"2A",X"01",X"FA",X"15",X"D0",X"BF",X"A8",X"F6",X"13",X"7D",X"25",X"A8",X"57",
		X"41",X"57",X"C0",X"FF",X"00",X"A9",X"0A",X"E0",X"BF",X"B4",X"FF",X"2A",X"75",X"5F",X"48",X"0A",
		X"2A",X"09",X"91",X"D2",X"AE",X"DA",X"DF",X"5A",X"8B",X"A8",X"00",X"35",X"51",X"8B",X"EE",X"AD",
		X"6F",X"D5",X"57",X"6D",X"81",X"94",X"2A",X"D0",X"7F",X"00",X"FB",X"05",X"E8",X"1B",X"80",X"BE",
		X"AA",X"FE",X"2F",X"F2",X"5F",X"D2",X"2B",X"00",X"70",X"01",X"F4",X"AB",X"F4",X"BF",X"A0",X"FF",
		X"02",X"F8",X"17",X"A0",X"2F",X"80",X"FF",X"02",X"F4",X"57",X"AA",X"4D",X"55",X"15",X"F0",X"F3",
		X"C1",X"17",X"80",X"FF",X"01",X"FC",X"02",X"C0",X"7F",X"D0",X"FF",X"BB",X"5A",X"5D",X"00",X"C0",
		X"36",X"00",X"7E",X"05",X"E8",X"5F",X"AB",X"FE",X"3A",X"40",X"5A",X"05",X"F0",X"FF",X"D1",X"57",
		X"93",X"42",X"FA",X"82",X"84",X"FF",X"00",X"F0",X"1F",X"F0",X"1F",X"00",X"F0",X"8F",X"BE",X"2A",
		X"5D",X"EA",X"D7",X"57",X"A5",X"B6",X"80",X"2B",X"78",X"25",X"A8",X"76",X"0A",X"FC",X"07",X"78",
		X"05",X"FB",X"03",X"E0",X"7F",X"80",X"FF",X"03",X"F0",X"7F",X"00",X"7C",X"05",X"AD",X"F6",X"03",
		X"D8",X"FF",X"40",X"57",X"00",X"F0",X"03",X"FE",X"5F",X"D4",X"F6",X"22",X"B5",X"2A",X"C0",X"2A",
		X"A5",X"FF",X"77",X"A9",X"05",X"5F",X"00",X"F8",X"03",X"00",X"FF",X"83",X"FE",X"07",X"D1",X"0F",
		X"80",X"FF",X"80",X"5F",X"2B",X"FA",X"1F",X"40",X"6A",X"05",X"C0",X"7F",X"E8",X"55",X"5D",X"F0",
		X"15",X"F0",X"4F",X"A8",X"AE",X"A0",X"FF",X"05",X"F8",X"3F",X"00",X"FF",X"0F",X"E0",X"0F",X"80",
		X"D6",X"0A",X"FC",X"5F",X"AA",X"AA",X"BF",X"90",X"00",X"80",X"4A",X"D0",X"FE",X"DF",X"FF",X"BF",
		X"2A",X"80",X"2F",X"00",X"3F",X"00",X"FE",X"03",X"FA",X"1F",X"C0",X"FF",X"81",X"AA",X"03",X"F0",
		X"87",X"FA",X"45",X"1F",X"C0",X"3F",X"E4",X"5F",X"09",X"F0",X"1F",X"80",X"7F",X"00",X"FD",X"1F",
		X"60",X"0F",X"40",X"D5",X"75",X"FB",X"1F",X"F4",X"2F",X"80",X"15",X"2A",X"88",X"74",X"E1",X"9F",
		X"E0",X"FF",X"0F",X"EA",X"0F",X"80",X"57",X"E0",X"DE",X"16",X"C0",X"0F",X"C0",X"AF",X"7F",X"E8",
		X"FF",X"01",X"FC",X"02",X"D8",X"03",X"00",X"17",X"80",X"FF",X"47",X"FF",X"4F",X"74",X"09",X"C0",
		X"FF",X"B5",X"0F",X"80",X"36",X"10",X"FD",X"05",X"EC",X"0F",X"F4",X"0F",X"E0",X"17",X"00",X"F7",
		X"0B",X"D0",X"FF",X"A3",X"3B",X"A9",X"03",X"E0",X"7F",X"00",X"FE",X"0F",X"F0",X"0F",X"00",X"7E",
		X"80",X"FE",X"57",X"F4",X"5F",X"C8",X"5F",X"00",X"DD",X"02",X"E0",X"3F",X"F0",X"2F",X"5D",X"A5",
		X"8A",X"E4",X"F2",X"EF",X"AA",X"24",X"40",X"0A",X"D0",X"2F",X"C0",X"BF",X"00",X"FA",X"1F",X"FC",
		X"7F",X"A9",X"40",X"BF",X"52",X"05",X"5D",X"00",X"7C",X"40",X"97",X"B6",X"55",X"AD",X"F2",X"15",
		X"F0",X"FF",X"4B",X"6A",X"07",X"00",X"FF",X"03",X"D0",X"55",X"D4",X"FE",X"5F",X"44",X"FA",X"03",
		X"92",X"00",X"50",X"25",X"DD",X"FE",X"6F",X"FB",X"7F",X"52",X"0D",X"00",X"02",X"E2",X"5B",X"D4",
		X"FE",X"05",X"91",X"7F",X"00",X"FE",X"3F",X"C0",X"FF",X"00",X"70",X"05",X"D1",X"7F",X"85",X"FF",
		X"47",X"6D",X"01",X"50",X"AB",X"AA",X"15",X"D0",X"3F",X"F4",X"4F",X"00",X"B0",X"16",X"B1",X"DF",
		X"FF",X"AB",X"FE",X"22",X"48",X"24",X"00",X"BE",X"00",X"FE",X"F7",X"7F",X"A5",X"AA",X"84",X"54",
		X"97",X"80",X"02",X"A8",X"45",X"AD",X"FC",X"AF",X"FA",X"DB",X"BF",X"00",X"68",X"05",X"00",X"FF",
		X"83",X"FA",X"07",X"D2",X"FE",X"03",X"EA",X"02",X"AA",X"DA",X"B7",X"F4",X"42",X"5D",X"89",X"24",
		X"15",X"D9",X"7F",X"D3",X"5F",X"A4",X"48",X"20",X"7C",X"05",X"E8",X"0D",X"A0",X"37",X"D1",X"FB",
		X"5F",X"F7",X"FF",X"01",X"FA",X"09",X"00",X"02",X"80",X"BD",X"DF",X"D5",X"3D",X"F5",X"5F",X"D4",
		X"16",X"00",X"56",X"11",X"49",X"D5",X"DE",X"D5",X"5E",X"69",X"AB",X"AD",X"6A",X"D5",X"2B",X"00",
		X"55",X"00",X"D0",X"6E",X"D5",X"46",X"F6",X"AF",X"FE",X"BF",X"80",X"FE",X"05",X"6A",X"01",X"00",
		X"36",X"D1",X"BF",X"A5",X"FE",X"1F",X"F9",X"2D",X"00",X"54",X"04",X"92",X"DA",X"8A",X"FE",X"7F",
		X"D5",X"AD",X"5A",X"D5",X"BE",X"2A",X"41",X"00",X"00",X"AA",X"24",X"EC",X"7F",X"F5",X"DF",X"D4",
		X"8A",X"B4",X"22",X"92",X"A8",X"AA",X"DF",X"55",X"FF",X"17",X"A9",X"15",X"00",X"D4",X"4A",X"F7",
		X"AA",X"24",X"7D",X"00",X"6E",X"08",X"41",X"FE",X"5F",X"FD",X"17",X"E8",X"5D",X"25",X"22",X"A5",
		X"BF",X"12",X"55",X"11",X"00",X"B5",X"A8",X"FF",X"82",X"FE",X"AF",X"2A",X"90",X"2A",X"52",X"25",
		X"FD",X"0B",X"F4",X"FF",X"0A",X"F5",X"17",X"40",X"2B",X"01",X"B6",X"93",X"94",X"6A",X"0B",X"ED",
		X"AF",X"FD",X"FA",X"1B",X"40",X"AF",X"00",X"B2",X"AA",X"B4",X"DD",X"1A",X"01",X"70",X"0B",X"E8",
		X"BF",X"20",X"FF",X"1F",X"FC",X"0F",X"A8",X"24",X"48",X"6D",X"01",X"FD",X"25",X"EA",X"AE",X"2A",
		X"6A",X"11",X"C9",X"FF",X"09",X"FE",X"03",X"E8",X"4A",X"6A",X"B7",X"A8",X"FF",X"04",X"3D",X"01",
		X"54",X"A5",X"4A",X"2B",X"A9",X"EA",X"DF",X"57",X"6A",X"95",X"5A",X"45",X"05",X"E8",X"15",X"F8",
		X"1F",X"A0",X"5F",X"01",X"ED",X"07",X"E0",X"9F",X"A8",X"FB",X"17",X"F4",X"BF",X"90",X"A4",X"04",
		X"80",X"37",X"48",X"77",X"BB",X"FD",X"57",X"EA",X"02",X"40",X"89",X"40",X"BA",X"AD",X"FE",X"FF",
		X"6D",X"A5",X"4A",X"90",X"04",X"AA",X"00",X"7D",X"4B",X"BB",X"2B",X"AA",X"FB",X"81",X"FE",X"4A",
		X"2A",X"A9",X"02",X"88",X"5A",X"4B",X"F8",X"FF",X"AA",X"AD",X"0A",X"80",X"77",X"11",X"52",X"5B",
		X"D2",X"FF",X"AD",X"5A",X"55",X"05",X"41",X"68",X"2B",X"A1",X"FF",X"4A",X"AA",X"BE",X"42",X"55",
		X"A2",X"0A",X"FA",X"9B",X"68",X"6B",X"15",X"FD",X"2B",X"E8",X"15",X"02",X"A9",X"0A",X"B4",X"57",
		X"FD",X"F7",X"7B",X"49",X"25",X"A5",X"08",X"84",X"90",X"90",X"BE",X"93",X"FA",X"2F",X"D5",X"BF",
		X"94",X"ED",X"0A",X"A8",X"04",X"74",X"5F",X"01",X"FD",X"09",X"B4",X"76",X"AD",X"5A",X"05",X"5D",
		X"A0",X"FE",X"11",X"DD",X"5B",X"40",X"7F",X"01",X"FC",X"26",X"C8",X"BE",X"89",X"FA",X"56",X"8A",
		X"B2",X"57",X"AA",X"56",X"81",X"A2",X"14",X"D4",X"7B",X"FD",X"5B",X"ED",X"56",X"52",X"6A",X"01",
		X"80",X"94",X"A4",X"DB",X"D5",X"FB",X"AB",X"FE",X"07",X"02",X"49",X"40",X"D2",X"26",X"D4",X"FE",
		X"A5",X"FE",X"BB",X"DA",X"BE",X"0A",X"A0",X"0A",X"C2",X"04",X"D0",X"B6",X"D5",X"F7",X"55",X"7D",
		X"AB",X"6C",X"15",X"B4",X"2B",X"EA",X"AD",X"00",X"E9",X"DB",X"AA",X"02",X"42",X"A9",X"6A",X"5F",
		X"49",X"55",X"ED",X"02",X"BA",X"02",X"B8",X"AB",X"FA",X"FF",X"56",X"B7",X"04",X"AA",X"54",X"ED",
		X"2A",X"80",X"0A",X"40",X"5F",X"A1",X"FE",X"56",X"BA",X"9F",X"C8",X"5D",X"15",X"88",X"AA",X"A4",
		X"7B",X"ED",X"BE",X"BB",X"02",X"55",X"00",X"6A",X"17",X"80",X"BE",X"22",X"7F",X"6B",X"BB",X"AD",
		X"92",X"2A",X"A5",X"4A",X"F5",X"55",X"52",X"DB",X"0A",X"D2",X"02",X"20",X"E9",X"16",X"F8",X"7F",
		X"AA",X"FF",X"25",X"B0",X"1F",X"A0",X"DA",X"22",X"95",X"0A",X"D2",X"AD",X"D4",X"BF",X"65",X"25",
		X"55",X"5F",X"C0",X"9F",X"38",X"A2",X"0F",X"BE",X"D0",X"6B",X"AA",X"C0",X"0F",X"F8",X"4A",X"BA",
		X"F5",X"02",X"AB",X"4A",X"D4",X"6E",X"69",X"55",X"A5",X"F2",X"8A",X"92",X"2E",X"FA",X"A2",X"2E",
		X"D2",X"52",X"17",X"6A",X"7D",X"89",X"FC",X"01",X"5B",X"85",X"FA",X"85",X"BE",X"A2",X"16",X"55",
		X"E8",X"A6",X"B4",X"6F",X"01",X"7D",X"64",X"E4",X"07",X"6A",X"57",X"49",X"7C",X"D1",X"15",X"FA",
		X"95",X"28",X"B5",X"82",X"FA",X"5A",X"ED",X"15",X"D0",X"D2",X"0B",X"DA",X"BE",X"54",X"D4",X"D2",
		X"05",X"FE",X"05",X"79",X"91",X"AA",X"EC",X"52",X"F5",X"A5",X"54",X"49",X"C5",X"56",X"AA",X"BD",
		X"52",X"A5",X"04",X"FE",X"0A",X"F9",X"41",X"5D",X"AA",X"BA",X"8A",X"D2",X"0E",X"AD",X"B4",X"9A",
		X"AA",X"EA",X"00",X"7F",X"05",X"FF",X"A8",X"E8",X"02",X"F6",X"85",X"BE",X"89",X"DA",X"0A",X"54",
		X"57",X"E8",X"2B",X"57",X"C1",X"4F",X"B0",X"07",X"F5",X"1D",X"D0",X"1B",X"BA",X"B0",X"57",X"A5",
		X"05",X"EA",X"07",X"FE",X"01",X"DF",X"14",X"72",X"4D",X"B5",X"A4",X"7E",X"E0",X"25",X"7C",X"0B",
		X"7A",X"45",X"EA",X"2B",X"68",X"5D",X"C1",X"9A",X"4E",X"F1",X"15",X"93",X"2D",X"15",X"DB",X"E0",
		X"1E",X"F2",X"2D",X"D4",X"C5",X"06",X"FC",X"49",X"A9",X"5F",X"A0",X"56",X"AA",X"E9",X"0B",X"57",
		X"BA",X"A0",X"55",X"BE",X"60",X"9F",X"22",X"F4",X"0B",X"FC",X"6A",X"A0",X"1F",X"28",X"F5",X"0B",
		X"FC",X"05",X"49",X"7F",X"C0",X"5F",X"02",X"FD",X"41",X"AA",X"2F",X"D0",X"4F",X"C8",X"3E",X"50",
		X"7B",X"05",X"FA",X"03",X"FA",X"AA",X"A0",X"3F",X"D0",X"57",X"41",X"FD",X"80",X"6F",X"15",X"F4",
		X"07",X"7C",X"55",X"D0",X"0F",X"D4",X"AF",X"40",X"BF",X"80",X"5F",X"21",X"FD",X"02",X"FD",X"82",
		X"F4",X"15",X"E4",X"2F",X"D0",X"B7",X"A0",X"BE",X"02",X"7B",X"85",X"FA",X"82",X"FA",X"44",X"7D",
		X"01",X"FD",X"09",X"EA",X"17",X"E8",X"17",X"E8",X"27",X"68",X"3F",X"A0",X"5F",X"A0",X"5F",X"81",
		X"7E",X"40",X"BF",X"A0",X"BD",X"90",X"BE",X"80",X"BF",X"40",X"BF",X"A0",X"AF",X"A0",X"5D",X"D4",
		X"55",X"D4",X"56",X"A9",X"92",X"6F",X"40",X"7F",X"A0",X"AF",X"D0",X"2E",X"E4",X"17",X"E8",X"0B",
		X"FA",X"81",X"7D",X"05",X"FD",X"02",X"BE",X"D0",X"16",X"7A",X"57",X"92",X"2F",X"D0",X"0B",X"FA",
		X"41",X"7D",X"05",X"7D",X"89",X"BA",X"D0",X"0F",X"EA",X"15",X"D4",X"15",X"F4",X"07",X"F5",X"85",
		X"DE",X"40",X"6D",X"45",X"3B",X"68",X"2F",X"74",X"AB",X"D4",X"0A",X"BD",X"40",X"FB",X"42",X"77",
		X"29",X"2F",X"D0",X"1D",X"F0",X"17",X"D4",X"07",X"F9",X"05",X"FA",X"45",X"B6",X"25",X"B5",X"80",
		X"3F",X"E0",X"5F",X"D0",X"57",X"E0",X"17",X"E8",X"8B",X"F4",X"12",X"BD",X"88",X"FE",X"80",X"7F",
		X"80",X"5F",X"C0",X"7E",X"D0",X"2B",X"E9",X"85",X"F4",X"05",X"FA",X"82",X"7E",X"81",X"7D",X"05",
		X"7D",X"A0",X"5F",X"A0",X"5F",X"C0",X"9F",X"E0",X"4B",X"7A",X"89",X"6E",X"A1",X"5E",X"81",X"BF",
		X"80",X"3F",X"C8",X"5E",X"51",X"2D",X"EA",X"05",X"BD",X"45",X"FA",X"0A",X"FA",X"22",X"56",X"75",
		X"81",X"7E",X"05",X"FD",X"05",X"BA",X"A5",X"A8",X"BE",X"40",X"FD",X"02",X"7B",X"A2",X"37",X"E8",
		X"15",X"DA",X"21",X"FD",X"40",X"3F",X"E0",X"0F",X"A9",X"0B",X"FD",X"04",X"FD",X"40",X"3F",X"E0",
		X"1F",X"F0",X"0B",X"FA",X"02",X"7B",X"A1",X"57",X"F4",X"02",X"FB",X"01",X"7F",X"C0",X"57",X"A8",
		X"17",X"7A",X"41",X"5F",X"C8",X"0F",X"F4",X"0B",X"FC",X"42",X"BE",X"A0",X"17",X"EA",X"03",X"FD",
		X"02",X"7F",X"C0",X"57",X"74",X"05",X"7F",X"C0",X"5F",X"D0",X"17",X"F4",X"09",X"9F",X"D0",X"17",
		X"E8",X"0F",X"F4",X"A2",X"2E",X"E8",X"17",X"F8",X"05",X"7B",X"C8",X"1E",X"E8",X"0B",X"79",X"91",
		X"5E",X"E8",X"0B",X"FC",X"01",X"7F",X"41",X"2F",X"F4",X"42",X"5F",X"D0",X"2E",X"A9",X"2B",X"B9",
		X"48",X"AF",X"E0",X"0F",X"F8",X"81",X"3E",X"F0",X"17",X"F8",X"41",X"BD",X"D0",X"07",X"FA",X"05",
		X"BD",X"A2",X"2B",X"F8",X"05",X"7E",X"81",X"1F",X"D4",X"0B",X"7E",X"A0",X"1F",X"F8",X"09",X"7E",
		X"41",X"5F",X"D0",X"07",X"7D",X"41",X"3F",X"D0",X"17",X"7C",X"81",X"5F",X"D0",X"07",X"FE",X"02",
		X"3F",X"D0",X"17",X"7A",X"91",X"7A",X"50",X"2F",X"F4",X"81",X"BE",X"D0",X"0B",X"FE",X"80",X"5F",
		X"E0",X"07",X"BE",X"D0",X"2E",X"F4",X"09",X"7D",X"E0",X"07",X"7D",X"C1",X"0F",X"FC",X"40",X"1F",
		X"F4",X"03",X"7D",X"41",X"2F",X"7A",X"A1",X"5E",X"D0",X"83",X"FA",X"82",X"7E",X"B0",X"A3",X"1E",
		X"E8",X"87",X"F4",X"05",X"7D",X"A0",X"2F",X"E8",X"83",X"BE",X"A0",X"1F",X"F0",X"05",X"BF",X"E0",
		X"0B",X"7D",X"41",X"2F",X"E8",X"83",X"BE",X"A0",X"1F",X"F8",X"03",X"7E",X"E0",X"07",X"FA",X"81",
		X"5F",X"D0",X"0B",X"7E",X"C0",X"9F",X"D0",X"43",X"BD",X"60",X"4F",X"F4",X"82",X"BD",X"A0",X"2E",
		X"EA",X"A2",X"5F",X"E0",X"0F",X"F4",X"42",X"5F",X"E0",X"17",X"F4",X"41",X"5F",X"F0",X"0B",X"7A",
		X"D0",X"4F",X"F0",X"03",X"3F",X"E4",X"0B",X"FA",X"C0",X"0F",X"F2",X"41",X"5F",X"E8",X"05",X"7D",
		X"C1",X"17",X"FA",X"C0",X"5E",X"F0",X"05",X"7D",X"D0",X"0F",X"7A",X"C1",X"0F",X"F8",X"83",X"3E",
		X"E8",X"0B",X"FC",X"A0",X"17",X"FA",X"40",X"5F",X"E8",X"05",X"3F",X"D0",X"0B",X"7D",X"E0",X"17",
		X"7C",X"C2",X"0F",X"FA",X"C0",X"0F",X"F8",X"05",X"7E",X"D0",X"07",X"7D",X"D0",X"07",X"FA",X"C0",
		X"17",X"7C",X"A1",X"0F",X"F4",X"03",X"AF",X"78",X"41",X"3F",X"E8",X"93",X"8E",X"F4",X"42",X"2F",
		X"F8",X"C1",X"0F",X"BC",X"A2",X"0E",X"7D",X"A0",X"0F",X"7A",X"C1",X"0F",X"7C",X"51",X"17",X"3E",
		X"C4",X"17",X"7A",X"C1",X"47",X"5E",X"E8",X"45",X"5D",X"D4",X"92",X"8D",X"F4",X"D0",X"17",X"7C",
		X"A1",X"0F",X"FA",X"C0",X"0F",X"7A",X"D0",X"17",X"7C",X"A1",X"0B",X"7D",X"D0",X"07",X"BD",X"F0",
		X"03",X"3F",X"F0",X"A1",X"5E",X"F0",X"05",X"1F",X"F4",X"A1",X"2E",X"F4",X"81",X"9F",X"F0",X"C8",
		X"27",X"F4",X"42",X"0F",X"7D",X"D0",X"07",X"7E",X"E0",X"07",X"7E",X"D0",X"07",X"7E",X"E0",X"07",
		X"7D",X"D0",X"0B",X"7E",X"D0",X"87",X"5E",X"E8",X"05",X"3F",X"D0",X"07",X"BD",X"D0",X"03",X"7F",
		X"E0",X"0B",X"3D",X"F2",X"41",X"9F",X"E0",X"0B",X"3D",X"D4",X"07",X"7D",X"D0",X"0B",X"FA",X"C1",
		X"17",X"F4",X"05",X"5F",X"F0",X"05",X"FD",X"C0",X"0F",X"7A",X"D0",X"07",X"FA",X"50",X"5F",X"E8",
		X"41",X"1F",X"F8",X"41",X"3B",X"E4",X"07",X"BD",X"E0",X"07",X"FC",X"42",X"2F",X"F4",X"0A",X"5F",
		X"B0",X"07",X"7D",X"A1",X"07",X"ED",X"83",X"5E",X"E8",X"03",X"5F",X"C1",X"0F",X"FC",X"82",X"17",
		X"7C",X"C1",X"1F",X"F0",X"83",X"5E",X"F0",X"03",X"7E",X"E0",X"17",X"7A",X"A1",X"07",X"7E",X"82",
		X"5F",X"F0",X"85",X"3E",X"F0",X"03",X"7D",X"D0",X"07",X"FD",X"C0",X"0F",X"BA",X"D0",X"17",X"FC",
		X"C0",X"2F",X"78",X"C1",X"0F",X"FC",X"82",X"1F",X"F8",X"81",X"2F",X"F8",X"05",X"6F",X"E8",X"02",
		X"3F",X"E8",X"85",X"3E",X"E8",X"85",X"1E",X"F8",X"0A",X"AF",X"F8",X"01",X"5F",X"F8",X"C0",X"17",
		X"7A",X"A4",X"87",X"7C",X"A8",X"8B",X"BC",X"E8",X"05",X"BF",X"E0",X"43",X"5F",X"F0",X"41",X"2F",
		X"F4",X"81",X"2F",X"F8",X"60",X"2F",X"F8",X"D0",X"07",X"FA",X"A0",X"0F",X"7E",X"E0",X"0B",X"7D",
		X"E0",X"83",X"3E",X"F0",X"03",X"1F",X"F4",X"C1",X"0F",X"7C",X"D1",X"03",X"7D",X"D1",X"45",X"2F",
		X"F8",X"82",X"8F",X"F8",X"C0",X"17",X"7C",X"A1",X"27",X"2E",X"F9",X"90",X"3E",X"F8",X"C0",X"0F",
		X"7E",X"E0",X"07",X"BD",X"D0",X"83",X"5E",X"F8",X"C0",X"17",X"7A",X"D0",X"0F",X"3A",X"F2",X"81",
		X"1F",X"F8",X"81",X"1F",X"FC",X"C0",X"0F",X"FC",X"42",X"27",X"3D",X"D1",X"55",X"87",X"BC",X"B0",
		X"07",X"BE",X"D0",X"85",X"3E",X"E8",X"89",X"17",X"7C",X"D0",X"07",X"3F",X"D0",X"0B",X"3D",X"F0",
		X"83",X"5E",X"F2",X"42",X"57",X"58",X"D3",X"B1",X"07",X"F9",X"A0",X"8F",X"F4",X"84",X"2F",X"F8",
		X"82",X"2F",X"2C",X"EB",X"18",X"DE",X"A4",X"A4",X"2F",X"F8",X"81",X"2F",X"F8",X"C2",X"07",X"FC",
		X"81",X"0F",X"7A",X"A1",X"0F",X"BE",X"E0",X"85",X"1F",X"F8",X"41",X"3F",X"F0",X"C1",X"17",X"F8",
		X"81",X"1F",X"F8",X"41",X"1F",X"7C",X"D0",X"0F",X"7C",X"A8",X"5B",X"F4",X"90",X"A7",X"E6",X"18",
		X"DA",X"C1",X"0F",X"F8",X"81",X"3F",X"F0",X"81",X"3E",X"F0",X"07",X"BE",X"D0",X"36",X"BC",X"81",
		X"5F",X"E0",X"0F",X"7C",X"E0",X"17",X"7A",X"A1",X"4F",X"E8",X"17",X"F4",X"02",X"BD",X"F0",X"03",
		X"7E",X"C1",X"2F",X"D8",X"81",X"BE",X"44",X"2F",X"F8",X"03",X"FE",X"80",X"3F",X"F0",X"21",X"3F",
		X"E8",X"43",X"EA",X"16",X"FA",X"88",X"17",X"EA",X"05",X"BF",X"80",X"1F",X"F4",X"81",X"BD",X"F0",
		X"85",X"7A",X"81",X"FE",X"C0",X"0F",X"FC",X"A0",X"1F",X"F0",X"03",X"FD",X"A0",X"2F",X"E8",X"43",
		X"3E",X"F0",X"0B",X"FA",X"82",X"2F",X"B4",X"A8",X"17",X"F8",X"05",X"BB",X"A2",X"47",X"7A",X"C8",
		X"4B",X"FA",X"86",X"BC",X"D0",X"07",X"7A",X"C2",X"0F",X"F8",X"81",X"3F",X"F0",X"41",X"1F",X"F4",
		X"05",X"5F",X"B0",X"07",X"5F",X"F0",X"05",X"5F",X"D0",X"0B",X"FA",X"41",X"1F",X"F4",X"C8",X"23",
		X"7C",X"41",X"3B",X"7E",X"E0",X"07",X"FC",X"A0",X"2F",X"B8",X"C3",X"17",X"BA",X"42",X"AF",X"2C",
		X"CE",X"E0",X"0B",X"EE",X"60",X"17",X"FA",X"81",X"1F",X"F8",X"C1",X"0F",X"F8",X"05",X"2F",X"F4",
		X"81",X"1F",X"F8",X"60",X"47",X"3B",X"E1",X"07",X"DD",X"D0",X"07",X"7D",X"E0",X"07",X"7E",X"E0",
		X"4B",X"2E",X"F4",X"82",X"2F",X"EA",X"A0",X"87",X"FE",X"A0",X"0B",X"1F",X"F8",X"41",X"17",X"FA",
		X"81",X"97",X"74",X"E4",X"27",X"3C",X"D2",X"31",X"9E",X"F4",X"10",X"9F",X"74",X"A8",X"47",X"78",
		X"CB",X"92",X"4E",X"E5",X"CA",X"86",X"1F",X"F0",X"07",X"3E",X"DA",X"A0",X"1F",X"E8",X"09",X"E7",
		X"36",X"B8",X"83",X"1E",X"FA",X"90",X"1E",X"76",X"E8",X"23",X"1D",X"F6",X"B0",X"86",X"65",X"AC",
		X"47",X"3C",X"D6",X"E2",X"0F",X"7E",X"50",X"C3",X"17",X"F8",X"C1",X"2B",X"7E",X"E0",X"07",X"6F",
		X"78",X"83",X"3E",X"F0",X"C1",X"0F",X"5E",X"F0",X"06",X"7D",X"E8",X"83",X"3F",X"B8",X"41",X"1F",
		X"E8",X"83",X"1E",X"BE",X"70",X"83",X"5F",X"B0",X"07",X"1F",X"F8",X"41",X"1F",X"F4",X"22",X"2F",
		X"F0",X"C1",X"87",X"F2",X"A2",X"07",X"7B",X"16",X"67",X"78",X"86",X"1D",X"7C",X"E8",X"83",X"BE",
		X"C0",X"0F",X"F8",X"83",X"0F",X"FC",X"C0",X"0F",X"FC",X"08",X"EB",X"70",X"D4",X"07",X"EA",X"17",
		X"3E",X"A8",X"63",X"FC",X"80",X"2F",X"A8",X"4F",X"3C",X"C9",X"4B",X"EC",X"0B",X"3E",X"E0",X"97",
		X"E8",X"C2",X"0F",X"7C",X"61",X"6A",X"19",X"FE",X"02",X"7E",X"E0",X"87",X"0E",X"7D",X"E8",X"47",
		X"3C",X"E0",X"3B",X"F8",X"C0",X"1E",X"E5",X"28",X"27",X"5F",X"05",X"F9",X"C0",X"BF",X"D0",X"27",
		X"B4",X"C7",X"09",X"47",X"39",X"5E",X"E1",X"2D",X"E8",X"08",X"EF",X"35",X"F4",X"88",X"CA",X"1F",
		X"F8",X"05",X"3E",X"A0",X"7F",X"01",X"7F",X"80",X"5F",X"A8",X"5F",X"D0",X"0B",X"EA",X"07",X"FE",
		X"80",X"DE",X"60",X"7D",X"A0",X"CE",X"41",X"7F",X"E0",X"07",X"FA",X"30",X"CE",X"43",X"8B",X"F1",
		X"05",X"FB",X"50",X"BA",X"15",X"FA",X"81",X"2F",X"A8",X"A7",X"A8",X"3E",X"F8",X"14",X"65",X"98",
		X"B7",X"41",X"2F",X"D0",X"1F",X"FC",X"C0",X"0F",X"F4",X"8B",X"D1",X"05",X"FB",X"88",X"5E",X"A2",
		X"37",X"D0",X"0D",X"6E",X"CB",X"06",X"FA",X"C1",X"2F",X"E8",X"81",X"3E",X"E8",X"0F",X"D4",X"07",
		X"7E",X"A0",X"3F",X"D0",X"0B",X"3B",X"AA",X"17",X"7A",X"C1",X"0E",X"FC",X"01",X"BF",X"E0",X"07",
		X"FC",X"81",X"3D",X"D8",X"A8",X"0F",X"DC",X"45",X"3D",X"D2",X"9A",X"1C",X"E5",X"0B",X"FC",X"40",
		X"5F",X"F8",X"81",X"2F",X"F0",X"43",X"2F",X"E8",X"07",X"BE",X"D0",X"85",X"AE",X"D0",X"2B",X"5E",
		X"C1",X"1F",X"F8",X"C0",X"0F",X"BE",X"E0",X"25",X"3D",X"E3",X"41",X"5E",X"F2",X"05",X"3F",X"E0",
		X"13",X"5F",X"F0",X"91",X"BA",X"B8",X"F0",X"07",X"F5",X"C0",X"0F",X"7A",X"A1",X"17",X"7A",X"85",
		X"6E",X"F8",X"82",X"96",X"5E",X"D0",X"07",X"BA",X"78",X"0B",X"7E",X"B0",X"32",X"C7",X"F8",X"80",
		X"5F",X"78",X"D5",X"E0",X"0F",X"F4",X"49",X"CB",X"74",X"C0",X"07",X"3F",X"87",X"31",X"1D",X"E1",
		X"03",X"AF",X"7A",X"5A",X"85",X"3A",X"EC",X"89",X"1E",X"F8",X"D0",X"47",X"79",X"C4",X"47",X"3C",
		X"E8",X"E3",X"05",X"FE",X"A0",X"1F",X"F0",X"F0",X"03",X"3F",X"F0",X"43",X"7C",X"D0",X"A1",X"0F",
		X"FE",X"20",X"C7",X"79",X"C2",X"07",X"BE",X"E8",X"95",X"16",X"F2",X"15",X"3E",X"E4",X"D8",X"8B",
		X"1E",X"F0",X"C3",X"71",X"83",X"53",X"7C",X"D0",X"43",X"1F",X"F4",X"11",X"CF",X"C1",X"1E",X"5E",
		X"F0",X"05",X"3F",X"F0",X"69",X"45",X"6B",X"C1",X"4F",X"F8",X"02",X"2F",X"7C",X"A0",X"1F",X"F8",
		X"41",X"AF",X"C3",X"A2",X"8B",X"78",X"07",X"3D",X"70",X"0F",X"FA",X"81",X"1F",X"F8",X"25",X"79",
		X"F0",X"05",X"7D",X"05",X"5F",X"F0",X"07",X"FC",X"C0",X"0F",X"FA",X"A0",X"2F",X"1C",X"97",X"70",
		X"4E",X"EA",X"03",X"BF",X"D0",X"9C",X"83",X"0F",X"F6",X"02",X"5F",X"C1",X"0F",X"BE",X"90",X"6E",
		X"E4",X"85",X"3C",X"D1",X"1F",X"F0",X"0B",X"FC",X"E0",X"C1",X"1F",X"D8",X"07",X"F4",X"13",X"5D",
		X"0B",X"F4",X"07",X"BE",X"A2",X"EA",X"05",X"BE",X"88",X"BE",X"24",X"F8",X"03",X"FE",X"A0",X"A6",
		X"2F",X"D4",X"43",X"95",X"FC",X"C0",X"17",X"A5",X"7D",X"81",X"6F",X"C1",X"0F",X"18",X"FD",X"82",
		X"CF",X"30",X"BA",X"03",X"D7",X"63",X"0D",X"36",X"A5",X"E9",X"03",X"FD",X"0A",X"FA",X"05",X"FC",
		X"03",X"7D",X"01",X"FF",X"80",X"BE",X"81",X"BE",X"44",X"7D",X"80",X"3F",X"A2",X"57",X"88",X"FD",
		X"C0",X"2F",X"E0",X"1F",X"C8",X"5B",X"D0",X"2F",X"D1",X"0B",X"EA",X"2D",X"F8",X"10",X"FD",X"82",
		X"3E",X"AC",X"CE",X"A2",X"6A",X"D1",X"07",X"E9",X"11",X"FD",X"81",X"0B",X"FB",X"02",X"DD",X"05",
		X"7E",X"C0",X"7D",X"E0",X"17",X"DC",X"21",X"7E",X"85",X"2B",X"51",X"77",X"38",X"EC",X"03",X"FE",
		X"02",X"5F",X"41",X"BF",X"84",X"53",X"FC",X"81",X"1F",X"E8",X"83",X"BE",X"A0",X"0F",X"EA",X"15",
		X"BC",X"A8",X"0B",X"F5",X"0A",X"5F",X"F0",X"03",X"3F",X"F0",X"27",X"E8",X"83",X"BE",X"E0",X"45",
		X"BE",X"C0",X"0F",X"FA",X"05",X"2F",X"FC",X"01",X"3F",X"E0",X"87",X"7A",X"A1",X"A5",X"7A",X"C8",
		X"07",X"F4",X"0B",X"2F",X"7C",X"48",X"5F",X"F0",X"06",X"AF",X"78",X"A8",X"0F",X"7E",X"01",X"1F",
		X"F9",X"A0",X"0F",X"7E",X"C0",X"17",X"FA",X"A4",X"07",X"7C",X"D1",X"4B",X"3A",X"A8",X"17",X"FA",
		X"A0",X"17",X"3D",X"C4",X"2B",X"7A",X"E8",X"03",X"7E",X"F0",X"86",X"3E",X"E0",X"07",X"7E",X"D0",
		X"8B",X"1E",X"F8",X"81",X"2F",X"7A",X"D0",X"17",X"F8",X"03",X"2F",X"7C",X"D0",X"0F",X"F8",X"A2",
		X"53",X"AE",X"E0",X"4B",X"4D",X"EA",X"40",X"3F",X"F0",X"0D",X"47",X"7D",X"A0",X"1F",X"F8",X"A0",
		X"5B",X"1E",X"E8",X"17",X"FC",X"C0",X"D1",X"07",X"FB",X"08",X"7E",X"E0",X"8B",X"0E",X"7D",X"E0",
		X"17",X"E8",X"0B",X"3E",X"F4",X"81",X"1F",X"F8",X"09",X"97",X"32",X"CB",X"2F",X"78",X"81",X"1F",
		X"FC",X"C0",X"17",X"7A",X"A1",X"17",X"74",X"8E",X"5E",X"E8",X"C2",X"3E",X"F4",X"21",X"1D",X"CE",
		X"03",X"3F",X"E0",X"BE",X"C0",X"0B",X"5E",X"8B",X"2F",X"F8",X"84",X"1F",X"F1",X"05",X"FD",X"40",
		X"5F",X"E0",X"33",X"3C",X"86",X"B7",X"F0",X"05",X"9D",X"31",X"FA",X"01",X"3F",X"F0",X"47",X"F8",
		X"20",X"1F",X"DA",X"F8",X"80",X"1F",X"EA",X"51",X"BC",X"95",X"78",X"0C",X"F9",X"03",X"F5",X"01",
		X"DF",X"03",X"7E",X"11",X"3F",X"41",X"5F",X"D4",X"3E",X"C0",X"F3",X"02",X"BF",X"01",X"5F",X"30",
		X"BF",X"02",X"7F",X"C0",X"9F",X"D0",X"25",X"25",X"7F",X"A0",X"0F",X"69",X"B5",X"D0",X"75",X"48",
		X"5F",X"01",X"7F",X"D0",X"3F",X"41",X"BE",X"80",X"BF",X"D4",X"82",X"0F",X"F4",X"17",X"6A",X"75",
		X"E0",X"2B",X"A2",X"5C",X"A5",X"5E",X"05",X"3E",X"55",X"ED",X"02",X"FE",X"02",X"7E",X"80",X"7F",
		X"C8",X"9B",X"80",X"7F",X"C2",X"3B",X"C0",X"5F",X"41",X"FB",X"80",X"7E",X"81",X"BE",X"05",X"FE",
		X"02",X"7E",X"0A",X"BB",X"07",X"EC",X"05",X"75",X"07",X"F4",X"07",X"EC",X"07",X"FC",X"0A",X"7A",
		X"8B",X"E8",X"07",X"DC",X"25",X"75",X"0B",X"F4",X"05",X"FD",X"85",X"D8",X"17",X"F4",X"03",X"7C",
		X"8B",X"7A",X"42",X"72",X"0D",X"3F",X"D0",X"07",X"DC",X"0F",X"7A",X"94",X"B3",X"4C",X"5E",X"D0",
		X"57",X"C8",X"0B",X"ED",X"0A",X"3F",X"E4",X"87",X"74",X"85",X"FC",X"02",X"7D",X"E0",X"1E",X"E8",
		X"13",X"FA",X"8A",X"2B",X"E3",X"82",X"7D",X"A1",X"07",X"F4",X"03",X"7F",X"E0",X"17",X"BA",X"05",
		X"7D",X"C8",X"2F",X"E0",X"87",X"FC",X"80",X"17",X"FA",X"A1",X"8F",X"D0",X"17",X"F9",X"82",X"2E",
		X"EA",X"05",X"7D",X"A0",X"1F",X"F8",X"81",X"3E",X"E8",X"03",X"BF",X"E0",X"03",X"BF",X"E0",X"0F",
		X"F8",X"05",X"BB",X"B4",X"41",X"5F",X"D0",X"17",X"BC",X"D0",X"17",X"7E",X"80",X"3F",X"F0",X"03",
		X"0F",X"FD",X"40",X"9F",X"E0",X"87",X"1E",X"7A",X"42",X"1F",X"FC",X"10",X"5F",X"78",X"C1",X"0F",
		X"FC",X"82",X"4F",X"E8",X"83",X"2F",X"BC",X"A0",X"1F",X"F8",X"82",X"2F",X"E8",X"C5",X"65",X"7C",
		X"A0",X"2F",X"E8",X"D1",X"13",X"FA",X"80",X"1F",X"79",X"45",X"17",X"7E",X"A0",X"2F",X"74",X"D4",
		X"07",X"FC",X"C0",X"AB",X"B4",X"D0",X"07",X"FE",X"40",X"0F",X"7D",X"E2",X"0B",X"FC",X"A0",X"17",
		X"7E",X"C0",X"0F",X"FC",X"81",X"0F",X"FA",X"C0",X"1F",X"F8",X"48",X"B7",X"B8",X"C0",X"17",X"F8",
		X"83",X"17",X"77",X"60",X"1F",X"E8",X"15",X"FA",X"D2",X"82",X"BD",X"A0",X"1F",X"68",X"87",X"F4",
		X"63",X"21",X"3F",X"E0",X"1F",X"F0",X"83",X"3E",X"D1",X"81",X"7E",X"E0",X"0F",X"F8",X"92",X"2E",
		X"EA",X"51",X"FA",X"02",X"7F",X"C0",X"1F",X"F8",X"81",X"3E",X"31",X"17",X"FC",X"B0",X"D6",X"52",
		X"BC",X"C2",X"35",X"42",X"3F",X"78",X"63",X"44",X"7F",X"50",X"0F",X"EC",X"91",X"FA",X"A0",X"5E",
		X"05",X"FD",X"82",X"7E",X"E0",X"5A",X"A1",X"2F",X"1D",X"E9",X"09",X"FC",X"05",X"FC",X"82",X"EE",
		X"29",X"B0",X"2F",X"D2",X"D6",X"02",X"FB",X"82",X"EA",X"0D",X"BA",X"2D",X"10",X"FE",X"C0",X"BF",
		X"40",X"7B",X"05",X"FD",X"40",X"3F",X"E0",X"0F",X"F4",X"27",X"C8",X"1D",X"E2",X"3F",X"A1",X"E8",
		X"05",X"BB",X"45",X"36",X"D5",X"D1",X"D0",X"8E",X"F8",X"0B",X"BA",X"C1",X"5B",X"72",X"A1",X"C2",
		X"FD",X"34",X"0B",X"F4",X"C1",X"5F",X"40",X"AF",X"92",X"7E",X"40",X"1F",X"75",X"51",X"55",X"D5",
		X"85",X"3F",X"B0",X"26",X"C3",X"DF",X"81",X"3C",X"85",X"5D",X"0B",X"F8",X"78",X"D4",X"91",X"B1",
		X"B4",X"07",X"BB",X"13",X"AA",X"7B",X"01",X"7E",X"C0",X"6F",X"A2",X"60",X"3F",X"C1",X"1F",X"C8",
		X"7E",X"C2",X"BA",X"40",X"DE",X"92",X"F3",X"2A",X"43",X"39",X"B4",X"FD",X"58",X"15",X"D4",X"87",
		X"58",X"0F",X"3F",X"D0",X"07",X"F8",X"03",X"EA",X"2F",X"E0",X"0F",X"E8",X"0F",X"AC",X"BD",X"80",
		X"7F",X"C0",X"2F",X"A8",X"5E",X"90",X"7B",X"41",X"7F",X"82",X"5F",X"C0",X"5F",X"50",X"5F",X"A0",
		X"57",X"D0",X"AF",X"E0",X"0B",X"EA",X"1B",X"7C",X"85",X"6C",X"0B",X"7D",X"F0",X"25",X"EA",X"05",
		X"7A",X"C2",X"17",X"EC",X"03",X"FE",X"01",X"BF",X"40",X"2F",X"B9",X"A5",X"D4",X"48",X"5F",X"41",
		X"3F",X"E0",X"0F",X"FA",X"03",X"6D",X"CA",X"91",X"B7",X"D0",X"97",X"B0",X"0B",X"EA",X"81",X"7F",
		X"60",X"0F",X"F5",X"A2",X"17",X"F0",X"07",X"EA",X"17",X"F8",X"88",X"1B",X"F4",X"42",X"5F",X"D0",
		X"07",X"7E",X"C1",X"8F",X"E8",X"03",X"7F",X"C0",X"2F",X"F0",X"0B",X"DE",X"42",X"8F",X"BA",X"D0",
		X"17",X"F8",X"81",X"3F",X"D0",X"07",X"FA",X"D0",X"13",X"75",X"A1",X"1F",X"F0",X"05",X"5F",X"F1",
		X"05",X"BE",X"B0",X"87",X"78",X"61",X"0F",X"F5",X"81",X"BE",X"C0",X"2F",X"74",X"85",X"3E",X"F4",
		X"03",X"7E",X"E0",X"0D",X"FA",X"60",X"5F",X"F0",X"03",X"2F",X"E9",X"92",X"AE",X"68",X"4F",X"F0",
		X"03",X"BE",X"24",X"2F",X"7D",X"C0",X"1F",X"E0",X"83",X"BE",X"70",X"A7",X"E8",X"03",X"7B",X"A8",
		X"2E",X"AA",X"2F",X"D0",X"1F",X"F8",X"60",X"1F",X"B2",X"07",X"FE",X"80",X"5D",X"E0",X"83",X"BE",
		X"48",X"3F",X"85",X"3E",X"F8",X"CC",X"83",X"3E",X"61",X"19",X"A3",X"47",X"1F",X"C1",X"17",X"EC",
		X"55",X"D0",X"1F",X"F0",X"1B",X"E0",X"0F",X"FC",X"84",X"EA",X"5D",X"E0",X"07",X"D4",X"0F",X"F8",
		X"17",X"E8",X"56",X"F0",X"17",X"E0",X"0F",X"D4",X"0F",X"EC",X"2B",X"A0",X"3F",X"50",X"7B",X"41",
		X"FD",X"09",X"F4",X"05",X"F6",X"52",X"EA",X"EA",X"02",X"B7",X"85",X"3E",X"7A",X"41",X"7A",X"D0",
		X"5B",X"0D",X"E5",X"21",X"FE",X"01",X"7F",X"01",X"7F",X"40",X"3F",X"14",X"FD",X"01",X"FB",X"04",
		X"6F",X"51",X"F5",X"48",X"57",X"19",X"ED",X"90",X"25",X"EB",X"A0",X"3D",X"6B",X"85",X"06",X"9D",
		X"7A",X"E0",X"5F",X"A5",X"96",X"70",X"9F",X"22",X"CF",X"70",X"91",X"BB",X"C8",X"07",X"2B",X"9A",
		X"A8",X"96",X"FA",X"05",X"2E",X"F1",X"0F",X"FA",X"40",X"3F",X"D4",X"15",X"BD",X"A0",X"07",X"F5",
		X"05",X"3B",X"A9",X"6A",X"78",X"E8",X"07",X"FE",X"50",X"5F",X"4C",X"4B",X"A2",X"A5",X"17",X"FC",
		X"40",X"6B",X"74",X"A5",X"4B",X"EA",X"11",X"FE",X"80",X"5F",X"A8",X"BA",X"A6",X"E8",X"0D",X"F0",
		X"03",X"7E",X"05",X"5F",X"37",X"E8",X"21",X"B6",X"B6",X"8A",X"F4",X"29",X"45",X"1B",X"D4",X"97",
		X"C4",X"A2",X"3F",X"E0",X"0F",X"FA",X"A3",X"05",X"F9",X"03",X"FD",X"42",X"F8",X"C0",X"0F",X"B4",
		X"2D",X"BA",X"D4",X"86",X"FA",X"03",X"FA",X"18",X"FE",X"21",X"7A",X"C5",X"81",X"56",X"6B",X"28",
		X"FF",X"00",X"BF",X"80",X"BF",X"24",X"F5",X"05",X"F4",X"83",X"B6",X"25",X"C9",X"6A",X"85",X"FE",
		X"40",X"5F",X"D0",X"DE",X"05",X"FA",X"07",X"FC",X"02",X"F4",X"0B",X"F8",X"13",X"F0",X"0B",X"F5",
		X"17",X"F0",X"95",X"F4",X"26",X"F8",X"0B",X"FA",X"01",X"F5",X"44",X"6D",X"49",X"5D",X"E8",X"0F",
		X"E8",X"17",X"68",X"1F",X"F8",X"16",X"FA",X"04",X"1F",X"E0",X"3D",X"D0",X"4F",X"D0",X"37",X"E8",
		X"07",X"BE",X"A2",X"6A",X"A5",X"43",X"3D",X"E1",X"7C",X"01",X"3F",X"60",X"7F",X"C0",X"0F",X"D4",
		X"8B",X"BA",X"D4",X"17",X"E8",X"0F",X"E8",X"43",X"F4",X"0B",X"FA",X"81",X"3D",X"E1",X"2D",X"F8",
		X"0A",X"7E",X"C1",X"2F",X"E0",X"3E",X"E8",X"1A",X"EC",X"42",X"BE",X"E0",X"8B",X"C8",X"3F",X"F0",
		X"05",X"F3",X"09",X"BF",X"C0",X"5F",X"A0",X"2F",X"68",X"2D",X"E9",X"05",X"3E",X"E1",X"1F",X"A0",
		X"5F",X"F0",X"07",X"F8",X"07",X"FC",X"01",X"3F",X"28",X"BF",X"40",X"5F",X"D0",X"3E",X"60",X"2F",
		X"F4",X"25",X"D4",X"F3",X"40",X"5F",X"A0",X"5F",X"A0",X"3F",X"F0",X"0B",X"F0",X"0F",X"E8",X"17",
		X"D8",X"17",X"B4",X"79",X"A1",X"2F",X"A1",X"36",X"68",X"77",X"21",X"7B",X"11",X"3F",X"D8",X"A2",
		X"BE",X"50",X"2F",X"60",X"6F",X"30",X"1F",X"F0",X"AE",X"F2",X"14",X"EA",X"09",X"95",X"B6",X"AB",
		X"76",X"E0",X"E4",X"55",X"0B",X"95",X"5E",X"A0",X"1F",X"F0",X"1F",X"E8",X"1A",X"C4",X"7D",X"C0",
		X"3F",X"D0",X"1E",X"AC",X"46",X"73",X"AD",X"E9",X"2A",X"58",X"83",X"7E",X"41",X"3F",X"42",X"FD",
		X"80",X"FE",X"02",X"EE",X"C1",X"AE",X"46",X"79",X"28",X"AE",X"86",X"AF",X"62",X"2D",X"B4",X"7C",
		X"93",X"FA",X"02",X"5C",X"07",X"FA",X"C3",X"D0",X"57",X"91",X"F6",X"25",X"F8",X"03",X"EA",X"A5",
		X"A0",X"BF",X"82",X"BF",X"A0",X"BE",X"50",X"E5",X"A2",X"09",X"2F",X"F4",X"54",X"C5",X"0D",X"7A",
		X"26",X"F4",X"17",X"EC",X"15",X"D4",X"0B",X"EA",X"5B",X"89",X"FA",X"84",X"4F",X"50",X"FA",X"16",
		X"9A",X"5E",X"E0",X"03",X"F6",X"4B",X"76",X"15",X"FC",X"02",X"F5",X"51",X"5A",X"17",X"E8",X"4F",
		X"A0",X"3F",X"A8",X"5E",X"A0",X"96",X"A5",X"B8",X"AB",X"56",X"A7",X"49",X"AD",X"A2",X"DE",X"68",
		X"23",X"E8",X"2D",X"9A",X"6E",X"C8",X"A5",X"68",X"AF",X"B8",X"2B",X"5E",X"05",X"BE",X"E0",X"9B",
		X"6A",X"07",X"E2",X"59",X"9C",X"4F",X"D8",X"4F",X"40",X"5F",X"41",X"5F",X"B0",X"D7",X"02",X"6F",
		X"34",X"0F",X"85",X"2E",X"F4",X"07",X"FC",X"03",X"BF",X"A0",X"5D",X"8A",X"9E",X"FA",X"00",X"DA",
		X"07",X"9B",X"3E",X"50",X"3F",X"C0",X"7F",X"80",X"3F",X"C1",X"1F",X"CC",X"07",X"FA",X"02",X"FE",
		X"50",X"B7",X"49",X"70",X"0F",X"F2",X"95",X"A0",X"3F",X"E0",X"1B",X"B4",X"AB",X"12",X"FA",X"16",
		X"EA",X"0B",X"D4",X"0F",X"F0",X"17",X"B4",X"9F",X"A0",X"5E",X"81",X"7E",X"81",X"7D",X"41",X"FA",
		X"03",X"ED",X"13",X"F8",X"25",X"E8",X"2F",X"E0",X"17",X"E8",X"2E",X"B0",X"AF",X"A0",X"3F",X"A0",
		X"AE",X"48",X"BF",X"44",X"7D",X"05",X"FD",X"82",X"F6",X"22",X"AD",X"02",X"F5",X"16",X"E9",X"0B",
		X"F4",X"03",X"ED",X"0F",X"F0",X"07",X"F8",X"55",X"E8",X"0F",X"F8",X"15",X"A4",X"5F",X"A0",X"FE",
		X"02",X"FA",X"02",X"FA",X"05",X"BD",X"64",X"A5",X"2F",X"F0",X"07",X"D5",X"9D",X"A0",X"3F",X"A0",
		X"2F",X"A4",X"E7",X"05",X"FC",X"15",X"F8",X"DA",X"82",X"FA",X"00",X"7F",X"01",X"3F",X"6A",X"D2",
		X"57",X"F0",X"0B",X"B7",X"50",X"4B",X"92",X"5F",X"A8",X"6B",X"11",X"D2",X"D7",X"2A",X"5D",X"6B",
		X"81",X"0E",X"B1",X"5F",X"F0",X"22",X"4D",X"CE",X"05",X"FE",X"03",X"7D",X"EA",X"82",X"3F",X"A0",
		X"2F",X"A4",X"55",X"A9",X"7A",X"01",X"1F",X"E1",X"5F",X"90",X"5E",X"85",X"FA",X"A2",X"BA",X"2A",
		X"C4",X"1F",X"54",X"3E",X"A4",X"E2",X"4B",X"D2",X"0F",X"DA",X"15",X"DA",X"2A",X"2D",X"EA",X"AB",
		X"80",X"7F",X"40",X"BF",X"14",X"EA",X"0F",X"F8",X"03",X"F4",X"47",X"A2",X"5E",X"A9",X"14",X"EA",
		X"BA",X"8E",X"61",X"E7",X"96",X"A8",X"3F",X"70",X"23",X"90",X"D7",X"0E",X"F2",X"A6",X"B8",X"AB",
		X"50",X"3D",X"D4",X"F1",X"2B",X"90",X"9B",X"C4",X"BE",X"80",X"FF",X"02",X"FC",X"07",X"F4",X"2D",
		X"70",X"0F",X"A6",X"67",X"A0",X"6B",X"44",X"D7",X"54",X"AE",X"8A",X"6D",X"30",X"7D",X"46",X"7F",
		X"01",X"7D",X"01",X"FF",X"02",X"FE",X"05",X"BA",X"13",X"F8",X"0B",X"F8",X"16",X"D8",X"AF",X"A0",
		X"6F",X"82",X"FA",X"40",X"5F",X"15",X"5E",X"43",X"DA",X"05",X"FD",X"12",X"FA",X"0B",X"7A",X"0B",
		X"F4",X"05",X"F2",X"16",X"EA",X"15",X"D4",X"52",X"95",X"5D",X"7D",X"15",X"A2",X"17",X"F1",X"72",
		X"92",X"D4",X"07",X"F9",X"0B",X"F4",X"0B",X"F5",X"8A",X"25",X"F9",X"42",X"7D",X"00",X"F7",X"82",
		X"FE",X"40",X"7B",X"08",X"BF",X"94",X"DE",X"92",X"F4",X"16",X"54",X"55",X"D6",X"2B",X"A0",X"0F",
		X"B8",X"47",X"59",X"BE",X"23",X"74",X"4B",X"AA",X"BD",X"54",X"1A",X"A9",X"FD",X"AE",X"00",X"AD",
		X"94",X"05",X"2F",X"FD",X"97",X"14",X"E5",X"83",X"E8",X"56",X"B1",X"2D",X"A0",X"7E",X"E8",X"22",
		X"7F",X"20",X"7E",X"81",X"5B",X"84",X"DF",X"02",X"FF",X"00",X"FD",X"AA",X"55",X"2D",X"82",X"FB",
		X"50",X"7A",X"89",X"DB",X"00",X"75",X"85",X"3E",X"FD",X"30",X"AE",X"D0",X"0F",X"F4",X"17",X"7C",
		X"81",X"96",X"FA",X"8A",X"7A",X"05",X"F4",X"00",X"FB",X"45",X"AF",X"B2",X"02",X"BF",X"A0",X"7F",
		X"B1",X"04",X"97",X"61",X"3D",X"D3",X"1E",X"EA",X"02",X"F8",X"23",X"F9",X"43",X"51",X"9F",X"A1",
		X"3E",X"E8",X"13",X"74",X"41",X"3F",X"D2",X"1F",X"E8",X"03",X"FC",X"52",X"A9",X"B7",X"00",X"AF",
		X"82",X"7B",X"AC",X"37",X"D0",X"17",X"E8",X"8B",X"E8",X"0F",X"46",X"95",X"52",X"AF",X"98",X"FC",
		X"10",X"7B",X"01",X"BF",X"A1",X"BE",X"83",X"5E",X"40",X"FF",X"90",X"D7",X"50",X"4D",X"49",X"26",
		X"1F",X"F8",X"1B",X"78",X"61",X"E5",X"46",X"2B",X"AE",X"2E",X"74",X"43",X"F9",X"52",X"5E",X"80",
		X"5F",X"C5",X"57",X"D4",X"AB",X"90",X"4A",X"B5",X"AA",X"52",X"48",X"9F",X"08",X"7F",X"A1",X"7F",
		X"81",X"FE",X"01",X"5C",X"45",X"FB",X"05",X"EA",X"45",X"BD",X"90",X"FE",X"82",X"3A",X"8A",X"F6",
		X"86",X"49",X"5A",X"D2",X"52",X"F1",X"55",X"3E",X"05",X"D9",X"57",X"D4",X"17",X"F4",X"0F",X"48",
		X"5A",X"52",X"55",X"FB",X"AE",X"2A",X"50",X"E9",X"78",X"49",X"DF",X"80",X"BF",X"04",X"6F",X"A1",
		X"7A",X"85",X"4A",X"CA",X"DB",X"35",X"94",X"55",X"AA",X"B7",X"42",X"7D",X"05",X"A6",X"49",X"BC",
		X"CE",X"2A",X"D6",X"15",X"70",X"97",X"F8",X"AE",X"94",X"46",X"E9",X"29",X"79",X"8B",X"B2",X"4A",
		X"F4",X"07",X"E8",X"7A",X"8E",X"E2",X"8B",X"F8",X"16",X"8A",X"6F",X"21",X"BE",X"86",X"AA",X"A3",
		X"A8",X"54",X"0B",X"F5",X"27",X"F4",X"42",X"B6",X"CA",X"B9",X"3C",X"F1",X"45",X"94",X"3F",X"A4",
		X"5D",X"A8",X"D8",X"91",X"C8",X"1B",X"89",X"EC",X"2A",X"F7",X"1A",X"D2",X"B7",X"24",X"6F",X"15",
		X"B4",X"8B",X"B2",X"4A",X"25",X"4B",X"B5",X"2D",X"68",X"1F",X"A0",X"6F",X"C8",X"57",X"88",X"FE",
		X"14",X"D4",X"2B",X"F5",X"65",X"61",X"1E",X"2D",X"A8",X"D6",X"6F",X"40",X"9D",X"E2",X"95",X"12",
		X"ED",X"1B",X"70",X"2F",X"A2",X"2B",X"D4",X"5B",X"C8",X"EA",X"CA",X"2B",X"88",X"BE",X"E2",X"BE",
		X"48",X"55",X"15",X"69",X"49",X"A8",X"5B",X"3F",X"80",X"BF",X"82",X"BF",X"A0",X"47",X"52",X"AA",
		X"DE",X"8A",X"A6",X"33",X"98",X"6A",X"AF",X"55",X"DB",X"8A",X"4B",X"40",X"DF",X"13",X"A2",X"AA",
		X"41",X"AA",X"F2",X"57",X"1A",X"9C",X"E2",X"A9",X"CE",X"57",X"07",X"F9",X"10",X"47",X"D8",X"5D",
		X"9A",X"A4",X"77",X"2A",X"29",X"BB",X"5F",X"80",X"56",X"A7",X"07",X"38",X"8F",X"13",X"F8",X"E3",
		X"58",X"C3",X"3D",X"8A",X"4B",X"D1",X"2F",X"78",X"35",X"84",X"FE",X"82",X"6B",X"84",X"2E",X"95",
		X"1E",X"E5",X"13",X"FE",X"50",X"B0",X"0F",X"F8",X"17",X"F4",X"16",X"D4",X"2B",X"C9",X"B5",X"53",
		X"BB",X"00",X"7D",X"11",X"55",X"EB",X"21",X"85",X"17",X"FC",X"45",X"BE",X"6D",X"09",X"7E",X"81",
		X"7D",X"01",X"3F",X"41",X"75",X"91",X"EA",X"93",X"6E",X"41",X"5A",X"53",X"7E",X"81",X"FF",X"00",
		X"7F",X"40",X"FF",X"00",X"BF",X"41",X"AC",X"53",X"BA",X"5B",X"B0",X"BA",X"40",X"FA",X"15",X"57",
		X"A9",X"56",X"15",X"94",X"6B",X"CB",X"2B",X"7C",X"2D",X"F0",X"02",X"CB",X"95",X"3D",X"35",X"FB",
		X"90",X"0F",X"40",X"7F",X"95",X"2B",X"00",X"DF",X"53",X"35",X"82",X"76",X"09",X"FF",X"5A",X"B4",
		X"07",X"E0",X"5F",X"C2",X"C3",X"D0",X"47",X"E1",X"45",X"6A",X"8D",X"ED",X"2F",X"C5",X"3E",X"18",
		X"BE",X"28",X"1D",X"2A",X"35",X"16",X"4D",X"59",X"0A",X"D6",X"FF",X"12",X"CB",X"F9",X"0E",X"46",
		X"29",X"9E",X"87",X"28",X"25",X"55",X"2B",X"8A",X"FF",X"25",X"AB",X"EA",X"3F",X"00",X"4F",X"C5",
		X"2F",X"01",X"D5",X"A8",X"B6",X"A1",X"68",X"FD",X"A3",X"E2",X"FA",X"6B",X"29",X"C0",X"F2",X"A9",
		X"54",X"28",X"AA",X"5A",X"35",X"90",X"FE",X"5B",X"38",X"FF",X"29",X"18",X"2A",X"7D",X"14",X"2A",
		X"1A",X"1E",X"2B",X"2E",X"0A",X"FF",X"0B",X"EA",X"BE",X"5E",X"26",X"90",X"3C",X"8F",X"4A",X"94",
		X"52",X"66",X"6B",X"40",X"FA",X"77",X"A3",X"EA",X"FD",X"14",X"24",X"52",X"BE",X"85",X"94",X"84",
		X"AD",X"25",X"4D",X"42",X"FB",X"5F",X"51",X"BC",X"FE",X"55",X"82",X"44",X"B5",X"BA",X"14",X"28",
		X"55",X"AD",X"23",X"A8",X"FE",X"ED",X"12",X"7C",X"7D",X"B5",X"14",X"A0",X"2E",X"9D",X"0A",X"4A",
		X"96",X"95",X"A3",X"E2",X"AF",X"81",X"EA",X"FB",X"77",X"01",X"D2",X"A5",X"EA",X"48",X"51",X"29",
		X"B5",X"D4",X"54",X"F4",X"03",X"FA",X"07",X"EA",X"FF",X"05",X"49",X"A9",X"56",X"53",X"91",X"44",
		X"55",X"AD",X"4A",X"A2",X"F6",X"EB",X"AB",X"A2",X"FB",X"3B",X"0C",X"51",X"AC",X"96",X"32",X"14",
		X"A6",X"9A",X"2A",X"85",X"DA",X"5F",X"D3",X"8A",X"EA",X"7F",X"0B",X"21",X"A9",X"55",X"92",X"8A",
		X"A2",X"58",X"D4",X"9A",X"54",X"1F",X"A0",X"5F",X"EF",X"FF",X"0A",X"60",X"73",X"9A",X"92",X"32",
		X"2A",X"55",X"29",X"AD",X"4A",X"DA",X"FF",X"12",X"D4",X"FB",X"7B",X"15",X"14",X"2D",X"0D",X"8B",
		X"8A",X"42",X"A5",X"AA",X"15",X"55",X"1B",X"DB",X"15",X"FE",X"DF",X"6B",X"40",X"5A",X"A9",X"2A",
		X"51",X"2A",X"4A",X"2A",X"57",X"43",X"B9",X"AE",X"EF",X"B1",X"FA",X"FB",X"3A",X"04",X"3C",X"0D",
		X"4D",X"09",X"96",X"86",X"AA",X"A5",X"42",X"75",X"F7",X"E9",X"34",X"FB",X"BB",X"97",X"00",X"55",
		X"A5",X"4A",X"09",X"51",X"51",X"79",X"AA",X"A0",X"5C",X"DF",X"AE",X"9A",X"EB",X"FD",X"1E",X"04",
		X"5A",X"8E",X"46",X"25",X"21",X"A3",X"65",X"D5",X"50",X"BA",X"BE",X"AE",X"56",X"AF",X"F7",X"75",
		X"09",X"50",X"4D",X"AA",X"12",X"44",X"25",X"AA",X"CB",X"42",X"C5",X"E5",X"EB",X"75",X"59",X"7B",
		X"5F",X"4F",X"09",X"A4",X"A3",X"4A",X"42",X"C9",X"A4",X"B4",X"B3",X"24",X"D4",X"FA",X"FA",X"A7",
		X"72",X"FB",X"DE",X"0D",X"41",X"5A",X"8A",X"2A",X"11",X"55",X"28",X"5D",X"95",X"0A",X"A5",X"AF",
		X"F5",X"B6",X"A4",X"F7",X"75",X"BD",X"04",X"38",X"86",X"A6",X"08",X"95",X"A2",X"D4",X"55",X"A9",
		X"44",X"F5",X"59",X"DF",X"D2",X"FC",X"BA",X"DF",X"0A",X"A8",X"4A",X"4A",X"45",X"42",X"25",X"25",
		X"A5",X"AB",X"45",X"A1",X"E9",X"EE",X"F5",X"B4",X"75",X"F5",X"BE",X"AE",X"10",X"18",X"97",X"29",
		X"0A",X"C5",X"52",X"55",X"CB",X"D2",X"2A",X"32",X"AD",X"FE",X"2E",X"A5",X"BF",X"B5",X"EE",X"92",
		X"10",X"52",X"2A",X"2C",X"24",X"1A",X"0B",X"4B",X"2B",X"97",X"87",X"44",X"A7",X"E7",X"BB",X"B2",
		X"F5",X"7C",X"75",X"3B",X"80",X"2C",X"0D",X"2B",X"46",X"45",X"95",X"A5",X"69",X"D5",X"55",X"A8",
		X"AC",X"78",X"BD",X"5E",X"56",X"AF",X"DE",X"D3",X"0A",X"C2",X"61",X"A9",X"42",X"D1",X"A8",X"B4",
		X"18",X"AD",X"AA",X"3A",X"0D",X"A5",X"AA",X"DE",X"57",X"D5",X"6D",X"F5",X"AE",X"47",X"40",X"2A",
		X"53",X"15",X"8A",X"45",X"31",X"AD",X"68",X"3A",X"56",X"2F",X"4A",X"8B",X"54",X"FF",X"56",X"35",
		X"B7",X"DD",X"4E",X"B7",X"00",X"AC",X"A5",X"A8",X"24",X"A9",X"94",X"AC",X"4A",X"AA",X"AA",X"D7",
		X"45",X"51",X"A5",X"B2",X"7F",X"AB",X"D5",X"6B",X"EB",X"FA",X"29",X"20",X"55",X"A9",X"2A",X"88",
		X"5A",X"92",X"56",X"89",X"AA",X"55",X"DD",X"AA",X"24",X"A1",X"EA",X"EA",X"7D",X"55",X"7D",X"5D",
		X"AE",X"2E",X"81",X"2A",X"45",X"55",X"A4",X"4A",X"51",X"55",X"49",X"D5",X"62",X"EF",X"D2",X"6A",
		X"28",X"A9",X"7A",X"BA",X"7E",X"2B",X"DD",X"57",X"97",X"8A",X"12",X"95",X"4A",X"52",X"0A",X"A3",
		X"49",X"A5",X"A2",X"52",X"CD",X"B1",X"6C",X"AD",X"A8",X"1A",X"92",X"76",X"5D",X"75",X"DF",X"AA",
		X"F6",X"B6",X"12",X"2A",X"85",X"26",X"45",X"45",X"A2",X"AA",X"94",X"AA",X"22",X"B5",X"2A",X"AD",
		X"1D",X"5D",X"17",X"55",X"15",X"D5",X"D7",X"6A",X"EB",X"7B",X"D5",X"BA",X"AA",X"AA",X"10",X"95",
		X"16",X"91",X"AA",X"84",X"AA",X"AA",X"AA",X"A2",X"D2",X"AA",X"D2",X"5A",X"AA",X"F7",X"6A",X"29",
		X"D5",X"59",X"BC",X"D7",X"B4",X"AE",X"D7",X"2D",X"85",X"D2",X"48",X"45",X"A9",X"4A",X"C2",X"32",
		X"A8",X"AA",X"A8",X"AC",X"A4",X"AA",X"2A",X"65",X"B5",X"AC",X"6E",X"A9",X"BA",X"AD",X"89",X"56",
		X"95",X"7A",X"AD",X"5F",X"55",X"5F",X"2B",X"94",X"16",X"49",X"2B",X"85",X"A5",X"82",X"D6",X"42",
		X"A9",X"45",X"D5",X"AA",X"AA",X"AA",X"AA",X"D6",X"A9",X"AA",X"A4",X"DA",X"3A",X"AA",X"B7",X"BA",
		X"44",X"7B",X"49",X"7D",X"55",X"5D",X"7D",X"55",X"A8",X"4A",X"A9",X"2A",X"A9",X"12",X"52",X"55",
		X"29",X"95",X"A2",X"5A",X"29",X"55",X"A9",X"6A",X"55",X"55",X"55",X"95",X"7E",X"25",X"B5",X"4A",
		X"95",X"0A",X"FD",X"8F",X"8A",X"57",X"D1",X"B5",X"D5",X"6A",X"B5",X"AA",X"A8",X"4A",X"51",X"55",
		X"95",X"48",X"A9",X"52",X"A9",X"54",X"AA",X"AA",X"B4",X"2A",X"55",X"55",X"5D",X"5F",X"45",X"AD",
		X"4A",X"7B",X"95",X"CA",X"52",X"B5",X"AA",X"52",X"55",X"41",X"FC",X"57",X"51",X"35",X"1D",X"DD",
		X"5E",X"AA",X"2A",X"55",X"15",X"95",X"96",X"4A",X"4A",X"95",X"92",X"4A",X"45",X"55",X"95",X"AA",
		X"AA",X"AA",X"AB",X"64",X"55",X"B5",X"55",X"A9",X"AA",X"AF",X"28",X"AD",X"D7",X"52",X"95",X"20",
		X"FA",X"2F",X"51",X"3A",X"9F",X"6A",X"5B",X"95",X"96",X"54",X"55",X"95",X"94",X"AA",X"4A",X"4A",
		X"25",X"A5",X"AA",X"4A",X"55",X"A5",X"5A",X"D5",X"AA",X"54",X"ED",X"AA",X"54",X"AD",X"68",X"ED",
		X"52",X"5A",X"55",X"55",X"55",X"55",X"A5",X"C0",X"F8",X"5D",X"A1",X"7A",X"59",X"7B",X"55",X"54",
		X"52",X"D5",X"AA",X"54",X"55",X"A8",X"5D",X"24",X"B5",X"52",X"6A",X"55",X"6A",X"95",X"6A",X"AB",
		X"54",X"B5",X"52",X"57",X"A5",X"6A",X"A5",X"AA",X"AA",X"6A",X"95",X"A8",X"AB",X"A2",X"D5",X"4A",
		X"55",X"55",X"A5",X"AB",X"A2",X"55",X"A5",X"56",X"A5",X"56",X"05",X"CB",X"AB",X"AA",X"82",X"FA",
		X"AB",X"AA",X"56",X"D2",X"EA",X"A2",X"6A",X"91",X"6A",X"A5",X"AA",X"2A",X"55",X"95",X"AA",X"AA",
		X"AA",X"5A",X"55",X"55",X"AD",X"56",X"95",X"B2",X"7E",X"AA",X"AE",X"A8",X"AA",X"AA",X"5A",X"95",
		X"AA",X"AA",X"5A",X"AA",X"AA",X"2A",X"4A",X"D7",X"2A",X"46",X"FB",X"5B",X"8A",X"56",X"A5",X"5A",
		X"15",X"AD",X"4A",X"AA",X"AA",X"AA",X"AA",X"54",X"55",X"55",X"D5",X"AA",X"AA",X"AA",X"AA",X"5A",
		X"95",X"AA",X"AA",X"BA",X"2A",X"55",X"55",X"55",X"AB",X"A4",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"A8",X"AA",X"AA",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"54",X"AD",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"1A",X"AA",X"57",X"55",X"2B",X"AA",X"5F",X"54",
		X"55",X"55",X"55",X"AA",X"5A",X"52",X"5B",X"51",X"5D",X"A4",X"5A",X"95",X"AA",X"AA",X"AA",X"55",
		X"55",X"95",X"5A",X"97",X"AA",X"AA",X"4A",X"AD",X"AA",X"AA",X"4A",X"D5",X"4B",X"55",X"AB",X"D0",
		X"56",X"51",X"B5",X"95",X"AA",X"95",X"54",X"AB",X"D4",X"2A",X"A9",X"AE",X"AA",X"AA",X"2A",X"6A",
		X"2D",X"55",X"AD",X"AA",X"AA",X"AA",X"2A",X"B5",X"2A",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"55",X"55",X"D5",
		X"AA",X"6A",X"55",X"D5",X"55",X"55",X"95",X"D0",X"B5",X"50",X"FD",X"22",X"B5",X"A3",X"D4",X"AA",
		X"A2",X"B5",X"8A",X"AE",X"52",X"5A",X"8B",X"6A",X"55",X"AA",X"AB",X"52",X"5A",X"A5",X"EA",X"AA",
		X"4A",X"D5",X"92",X"DA",X"55",X"B1",X"2A",X"AA",X"AB",X"92",X"AA",X"AB",X"54",X"AB",X"A2",X"6A",
		X"55",X"55",X"55",X"55",X"95",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"B5",
		X"AA",X"AA",X"54",X"B5",X"AA",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"55",X"B5",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"92",X"AA",X"55",X"55",X"AD",X"AA",X"AA",X"EA",X"56",
		X"A2",X"AA",X"AA",X"AB",X"AA",X"AA",X"52",X"B5",X"AA",X"AA",X"AA",X"AA",X"AA",X"52",X"55",X"55",
		X"55",X"A5",X"AA",X"AA",X"AA",X"AA",X"D5",X"55",X"A9",X"AA",X"54",X"6D",X"A9",X"54",X"55",X"55",
		X"A9",X"AA",X"AA",X"54",X"55",X"51",X"55",X"B5",X"68",X"5D",X"D4",X"B6",X"88",X"AE",X"AA",X"5A",
		X"5D",X"5D",X"A0",X"E8",X"03",X"1A",X"B5",X"EA",X"82",X"A2",X"4E",X"FD",X"74",X"FB",X"23",X"AD",
		X"2E",X"20",X"00",X"48",X"45",X"ED",X"FE",X"FF",X"AD",X"92",X"12",X"7A",X"11",X"21",X"09",X"DA",
		X"52",X"FB",X"7F",X"AB",X"4A",X"42",X"AD",X"BA",X"B5",X"4A",X"55",X"2F",X"80",X"D4",X"4A",X"25",
		X"12",X"BD",X"77",X"A1",X"AB",X"4B",X"54",X"48",X"E8",X"4A",X"AB",X"6E",X"BB",X"F6",X"ED",X"92",
		X"6E",X"AD",X"44",X"95",X"EA",X"55",X"95",X"54",X"BD",X"82",X"4A",X"12",X"52",X"55",X"90",X"A2",
		X"86",X"54",X"A9",X"54",X"A5",X"2A",X"54",X"A9",X"EB",X"FF",X"6F",X"DB",X"EF",X"AA",X"AA",X"4A",
		X"B5",X"AA",X"AA",X"24",X"55",X"29",X"52",X"AA",X"90",X"10",X"10",X"89",X"4A",X"92",X"F6",X"6E",
		X"6F",X"6B",X"57",X"B5",X"ED",X"AD",X"BA",X"75",X"D5",X"5A",X"D5",X"DF",X"55",X"0B",X"AA",X"4A",
		X"04",X"42",X"48",X"42",X"88",X"AA",X"6A",X"6D",X"6B",X"55",X"A8",X"5E",X"D5",X"AD",X"E2",X"EE",
		X"D6",X"DE",X"FD",X"AE",X"AA",X"52",X"55",X"55",X"49",X"4A",X"22",X"25",X"AA",X"56",X"45",X"55",
		X"52",X"22",X"88",X"A4",X"D6",X"FA",X"6A",X"DD",X"76",X"55",X"55",X"45",X"95",X"94",X"AA",X"6A",
		X"D5",X"AB",X"56",X"44",X"54",X"AB",X"4A",X"AD",X"AA",X"5A",X"55",X"A5",X"FA",X"15",X"00",X"D5",
		X"55",X"95",X"7E",X"B5",X"B7",X"82",X"BA",X"5D",X"6D",X"15",X"A0",X"F6",X"AB",X"82",X"C2",X"FF",
		X"1F",X"00",X"80",X"FF",X"AF",X"96",X"E6",X"FF",X"00",X"00",X"C0",X"FF",X"47",X"40",X"FD",X"7F",
		X"21",X"B2",X"94",X"AA",X"2E",X"02",X"A8",X"FF",X"4A",X"D4",X"FF",X"6F",X"95",X"AA",X"D6",X"AD",
		X"0A",X"41",X"AA",X"44",X"00",X"48",X"A5",X"DA",X"AA",X"FA",X"FD",X"DB",X"A5",X"4A",X"55",X"49",
		X"A2",X"EA",X"FB",X"56",X"82",X"EA",X"52",X"48",X"48",X"F5",X"56",X"04",X"00",X"F8",X"7F",X"09",
		X"50",X"B4",X"6F",X"2F",X"3D",X"7F",X"4A",X"A4",X"46",X"BD",X"FF",X"12",X"48",X"DB",X"26",X"AA",
		X"FA",X"55",X"21",X"12",X"01",X"A4",X"42",X"80",X"D4",X"BA",X"A9",X"ED",X"FE",X"7F",X"7F",X"F7",
		X"AE",X"54",X"52",X"01",X"01",X"20",X"52",X"7F",X"BD",X"52",X"5B",X"FD",X"40",X"01",X"A8",X"B4",
		X"80",X"6E",X"FD",X"ED",X"FF",X"AB",X"2A",X"81",X"3F",X"00",X"00",X"FA",X"FF",X"FD",X"65",X"97",
		X"5E",X"00",X"00",X"F0",X"FF",X"C1",X"87",X"FE",X"FF",X"57",X"02",X"50",X"C0",X"0D",X"00",X"88",
		X"F4",X"8F",X"FA",X"AA",X"FA",X"27",X"AD",X"02",X"AD",X"AE",X"FC",X"01",X"00",X"F8",X"BB",X"A4",
		X"6F",X"DB",X"BF",X"22",X"00",X"F8",X"1F",X"00",X"D8",X"FF",X"FF",X"AE",X"5A",X"C8",X"16",X"49",
		X"E0",X"BF",X"00",X"50",X"89",X"1F",X"00",X"00",X"F8",X"FF",X"FF",X"BF",X"DF",X"05",X"00",X"C0",
		X"FF",X"AF",X"A8",X"FF",X"7F",X"01",X"80",X"56",X"00",X"00",X"40",X"FF",X"87",X"0A",X"58",X"FD",
		X"83",X"02",X"BC",X"BF",X"F4",X"A3",X"DF",X"3F",X"39",X"00",X"40",X"2D",X"DD",X"E8",X"FF",X"FF",
		X"7F",X"00",X"00",X"20",X"0B",X"A0",X"F5",X"DF",X"07",X"C0",X"1E",X"58",X"F8",X"03",X"00",X"F0",
		X"FC",X"FF",X"CB",X"2F",X"10",X"01",X"A8",X"D4",X"FF",X"FF",X"FE",X"97",X"00",X"00",X"F8",X"FD",
		X"03",X"00",X"3C",X"F8",X"E0",X"83",X"FF",X"FF",X"10",X"00",X"F4",X"07",X"27",X"FF",X"7A",X"01",
		X"00",X"D1",X"BF",X"8F",X"FC",X"FF",X"11",X"08",X"80",X"FB",X"D7",X"2F",X"24",X"A9",X"82",X"D6",
		X"FE",X"B7",X"10",X"49",X"01",X"3F",X"00",X"C0",X"E1",X"FF",X"FF",X"7F",X"FF",X"0B",X"10",X"80",
		X"FF",X"FF",X"C0",X"FF",X"AF",X"00",X"C0",X"2F",X"3F",X"08",X"F0",X"F7",X"07",X"2B",X"15",X"FE",
		X"5D",X"40",X"C9",X"FE",X"0B",X"00",X"1F",X"5D",X"00",X"80",X"FF",X"FF",X"DD",X"FF",X"D6",X"92",
		X"C0",X"0F",X"3D",X"FE",X"00",X"02",X"5C",X"F5",X"AB",X"06",X"80",X"54",X"01",X"F4",X"FF",X"FF",
		X"3F",X"60",X"00",X"00",X"F8",X"FF",X"05",X"E0",X"FC",X"8F",X"1F",X"5C",X"FE",X"7F",X"04",X"00",
		X"FE",X"1F",X"80",X"AE",X"BF",X"11",X"00",X"90",X"FE",X"0B",X"80",X"FA",X"D3",X"02",X"00",X"F0",
		X"FF",X"1F",X"E0",X"FF",X"3F",X"FC",X"01",X"06",X"3E",X"08",X"C0",X"FF",X"A1",X"DB",X"0B",X"00",
		X"F0",X"C3",X"BB",X"FF",X"43",X"00",X"20",X"FB",X"EB",X"04",X"FC",X"3F",X"00",X"E8",X"EB",X"FE",
		X"2F",X"FF",X"01",X"00",X"10",X"7F",X"FF",X"6F",X"E5",X"27",X"00",X"00",X"80",X"FF",X"7F",X"A5",
		X"44",X"FD",X"0A",X"80",X"5F",X"40",X"BF",X"02",X"C0",X"FF",X"17",X"00",X"FE",X"FF",X"07",X"B0",
		X"7F",X"A9",X"05",X"80",X"AF",X"5A",X"03",X"00",X"FE",X"BF",X"00",X"41",X"FF",X"FF",X"47",X"00",
		X"FB",X"2F",X"00",X"A0",X"FF",X"23",X"00",X"40",X"37",X"BD",X"55",X"A1",X"FF",X"FF",X"0A",X"E8",
		X"FF",X"03",X"90",X"92",X"BE",X"08",X"F8",X"51",X"09",X"14",X"F0",X"FF",X"17",X"55",X"55",X"05",
		X"00",X"C0",X"FF",X"FF",X"AF",X"12",X"E8",X"07",X"82",X"54",X"FF",X"11",X"54",X"42",X"F4",X"7F",
		X"00",X"ED",X"FF",X"75",X"01",X"E0",X"FF",X"5F",X"02",X"D0",X"FF",X"01",X"00",X"F8",X"2B",X"01",
		X"00",X"FD",X"F3",X"BB",X"07",X"6C",X"FD",X"52",X"C9",X"FF",X"AB",X"54",X"FA",X"5F",X"01",X"94",
		X"00",X"44",X"15",X"28",X"F5",X"4F",X"5F",X"15",X"92",X"00",X"C0",X"BD",X"E5",X"FF",X"67",X"FF",
		X"0B",X"12",X"00",X"F0",X"F7",X"DA",X"12",X"DD",X"FF",X"01",X"A0",X"02",X"40",X"5D",X"D5",X"7F",
		X"FA",X"F7",X"00",X"FD",X"03",X"00",X"28",X"5A",X"D1",X"AB",X"FF",X"AD",X"7D",X"7B",X"C9",X"15",
		X"00",X"F4",X"D5",X"BE",X"05",X"DA",X"4B",X"50",X"95",X"08",X"EA",X"D2",X"57",X"00",X"F4",X"7F",
		X"81",X"FA",X"FB",X"4F",X"14",X"22",X"80",X"DF",X"92",X"F6",X"25",X"2A",X"C0",X"6A",X"81",X"FE",
		X"7F",X"49",X"A4",X"08",X"ED",X"7F",X"55",X"55",X"3F",X"00",X"50",X"09",X"A2",X"DA",X"92",X"C8",
		X"FF",X"FF",X"55",X"AB",X"2A",X"21",X"01",X"50",X"FF",X"6E",X"A5",X"5A",X"55",X"24",X"29",X"95",
		X"44",X"FD",X"57",X"EF",X"BE",X"5D",X"84",X"F4",X"17",X"00",X"00",X"B0",X"55",X"81",X"FE",X"FF",
		X"42",X"A4",X"EA",X"FF",X"95",X"5A",X"69",X"F7",X"17",X"E8",X"56",X"00",X"95",X"04",X"60",X"B7",
		X"0A",X"94",X"FE",X"F7",X"EF",X"1F",X"00",X"A0",X"44",X"20",X"75",X"FF",X"DF",X"B5",X"D2",X"F7",
		X"95",X"5A",X"B5",X"00",X"80",X"04",X"00",X"60",X"7F",X"5F",X"F7",X"6D",X"AB",X"B5",X"54",X"F5",
		X"FF",X"0A",X"00",X"20",X"48",X"04",X"40",X"BA",X"B7",X"12",X"C8",X"FF",X"FF",X"FF",X"DD",X"EE",
		X"4B",X"00",X"04",X"A9",X"52",X"90",X"88",X"AA",X"7F",X"01",X"00",X"DD",X"BD",X"AD",X"FF",X"BB",
		X"65",X"4B",X"80",X"48",X"55",X"AB",X"2A",X"75",X"DB",X"5F",X"09",X"20",X"55",X"11",X"F7",X"6F",
		X"F5",X"6F",X"01",X"80",X"64",X"ED",X"0B",X"48",X"55",X"AB",X"2E",X"20",X"55",X"DF",X"55",X"50",
		X"FD",X"6F",X"DB",X"FD",X"DF",X"EA",X"2F",X"00",X"00",X"EA",X"FF",X"55",X"05",X"00",X"48",X"22",
		X"92",X"FE",X"7F",X"6F",X"53",X"FF",X"D5",X"4A",X"00",X"00",X"F4",X"FF",X"23",X"F4",X"B6",X"02",
		X"40",X"BA",X"B5",X"A4",X"12",X"F5",X"FF",X"2F",X"AA",X"AA",X"57",X"02",X"92",X"A4",X"5A",X"01",
		X"48",X"BB",X"2D",X"49",X"A8",X"FE",X"AB",X"76",X"5B",X"FF",X"15",X"04",X"D5",X"EE",X"96",X"48",
		X"84",X"AA",X"2A",X"91",X"2A",X"01",X"D4",X"6A",X"FB",X"FF",X"DB",X"04",X"F5",X"4F",X"90",X"50",
		X"84",X"56",X"BF",X"6D",X"6D",X"0D",X"20",X"29",X"05",X"50",X"DF",X"FF",X"24",X"25",X"81",X"1A",
		X"F0",X"3F",X"10",X"FA",X"E0",X"FF",X"FF",X"07",X"00",X"14",X"29",X"C8",X"AD",X"7E",X"BF",X"01",
		X"AF",X"EA",X"7F",X"13",X"01",X"48",X"7A",X"45",X"02",X"0A",X"A4",X"FB",X"B6",X"AF",X"FE",X"EF",
		X"D5",X"6F",X"90",X"0A",X"00",X"90",X"92",X"55",X"22",X"55",X"12",X"69",X"FF",X"F7",X"5F",X"AB",
		X"FB",X"D7",X"AE",X"04",X"24",X"00",X"A0",X"D4",X"B6",X"AB",X"24",X"69",X"5B",X"DB",X"B5",X"D4",
		X"05",X"F5",X"AE",X"F4",X"17",X"00",X"A1",X"FE",X"5B",X"A5",X"AA",X"6A",X"AB",X"02",X"91",X"FA",
		X"2B",X"D2",X"05",X"FE",X"03",X"00",X"28",X"FD",X"FF",X"5F",X"00",X"D2",X"8D",X"20",X"FA",X"FF",
		X"3F",X"00",X"60",X"DB",X"BE",X"49",X"54",X"25",X"09",X"24",X"A9",X"FF",X"AA",X"6A",X"6D",X"FD",
		X"82",X"A4",X"BA",X"FF",X"16",X"40",X"02",X"24",X"21",X"40",X"A5",X"FB",X"6F",X"F5",X"BF",X"6F",
		X"6B",X"A9",X"5A",X"B5",X"52",X"02",X"51",X"5A",X"00",X"02",X"D2",X"BD",X"57",X"AD",X"52",X"DD",
		X"56",X"48",X"D2",X"F6",X"96",X"00",X"00",X"AA",X"FF",X"FF",X"92",X"AA",X"FE",X"AB",X"6A",X"DB",
		X"5A",X"02",X"A0",X"56",X"2A",X"01",X"90",X"AA",X"A4",X"55",X"A9",X"5F",X"00",X"FE",X"0F",X"04",
		X"10",X"FE",X"7F",X"FF",X"01",X"FE",X"07",X"00",X"C0",X"FF",X"7F",X"90",X"60",X"77",X"5F",X"00",
		X"D5",X"DD",X"24",X"00",X"40",X"FF",X"96",X"08",X"FA",X"FF",X"47",X"AA",X"FA",X"FF",X"07",X"28",
		X"40",X"5B",X"00",X"40",X"E9",X"FF",X"02",X"50",X"FD",X"FF",X"55",X"B5",X"7D",X"2F",X"44",X"64",
		X"AB",X"0D",X"00",X"00",X"B5",X"ED",X"84",X"54",X"FF",X"F5",X"4A",X"94",X"6F",X"ED",X"2E",X"EA",
		X"5E",X"49",X"29",X"D0",X"BF",X"B4",X"52",X"A5",X"BF",X"DA",X"AB",X"00",X"58",X"00",X"AB",X"92",
		X"AA",X"92",X"7A",X"00",X"68",X"6D",X"97",X"FE",X"07",X"50",X"FE",X"FD",X"FF",X"BD",X"82",X"0A",
		X"01",X"C8",X"F6",X"FF",X"2D",X"90",X"40",X"52",X"49",X"54",X"AB",X"AE",X"40",X"80",X"D4",X"7E",
		X"D5",X"EE",X"FF",X"AF",X"50",X"B5",X"FF",X"77",X"05",X"20",X"20",X"25",X"41",X"EA",X"B6",X"57",
		X"91",X"AA",X"DD",X"DF",X"AA",X"54",X"AB",X"10",X"20",X"B5",X"BF",X"8A",X"08",X"40",X"6D",X"AB",
		X"D4",X"4A",X"7D",X"45",X"7F",X"6F",X"EF",X"6D",X"49",X"55",X"55",X"11",X"91",X"ED",X"AF",X"2A",
		X"88",X"D4",X"56",X"92",X"88",X"A4",X"54",X"55",X"AB",X"AA",X"7A",X"05",X"49",X"6A",X"F5",X"17",
		X"EA",X"AA",X"BB",X"5B",X"ED",X"DD",X"56",X"55",X"A0",X"44",X"AA",X"AA",X"2A",X"A2",X"42",X"FD",
		X"1F",X"00",X"40",X"FF",X"AF",X"D2",X"02",X"58",X"05",X"90",X"FA",X"FF",X"7F",X"42",X"51",X"FF",
		X"AF",X"AA",X"AA",X"94",X"00",X"00",X"AA",X"ED",X"12",X"48",X"ED",X"DF",X"12",X"B5",X"FF",X"DF",
		X"8A",X"40",X"49",X"AA",X"04",X"A4",X"05",X"91",X"84",X"F4",X"BF",X"DB",X"6A",X"FB",X"BF",X"4A",
		X"55",X"F7",X"6E",X"22",X"80",X"94",X"52",X"00",X"6A",X"EF",X"9A",X"10",X"D4",X"FD",X"B6",X"4A",
		X"F2",X"DE",X"0A",X"52",X"75",X"BF",X"AD",X"AA",X"A5",X"6D",X"15",X"A8",X"2D",X"A9",X"12",X"22",
		X"85",X"28",X"01",X"90",X"DE",X"AA",X"B7",X"F6",X"5F",X"55",X"D5",X"AA",X"F6",X"AA",X"56",X"BB",
		X"92",X"04",X"D5",X"AA",X"54",X"BF",X"40",X"42",X"24",X"75",X"EF",X"9A",X"10",X"25",X"89",X"A8",
		X"54",X"F7",X"DB",X"A5",X"7A",X"EF",X"5E",X"F5",X"FF",X"01",X"88",X"54",X"7D",X"6D",X"15",X"40",
		X"02",X"00",X"A4",X"FF",X"BF",X"AA",X"AA",X"6A",X"77",X"6B",X"ED",X"56",X"15",X"00",X"52",X"A2",
		X"AA",X"88",X"FA",X"7B",X"AB",X"A0",X"FE",X"FF",X"AB",X"14",X"55",X"12",X"10",X"A0",X"EE",X"AE",
		X"08",X"90",X"6C",X"77",X"57",X"FB",X"DF",X"4A",X"80",X"DA",X"EF",X"95",X"12",X"94",X"2A",X"42",
		X"68",X"FB",X"6E",X"03",X"A4",X"DA",X"AE",X"B5",X"A4",X"AA",X"94",X"52",X"49",X"7D",X"BF",X"D5",
		X"AA",X"A4",X"0A",X"A2",X"77",X"6B",X"B7",X"88",X"0A",X"44",X"55",X"49",X"55",X"55",X"FB",X"AA",
		X"AA",X"52",X"FF",X"AE",X"AA",X"2A",X"EA",X"5B",X"25",X"08",X"A9",X"2A",X"12",X"89",X"EA",X"7D",
		X"77",X"5B",X"BB",X"95",X"40",X"AA",X"9D",X"12",X"00",X"50",X"55",X"55",X"55",X"55",X"AB",X"AA",
		X"F7",X"FB",X"FF",X"B7",X"2A",X"49",X"92",X"54",X"55",X"49",X"04",X"02",X"94",X"AA",X"5A",X"D5",
		X"EE",X"56",X"55",X"FD",X"EF",X"6B",X"95",X"00",X"A9",X"94",X"A4",X"DA",X"6E",X"95",X"A4",X"D6",
		X"DE",X"96",X"A0",X"F6",X"EE",X"55",X"A5",X"94",X"92",X"10",X"22",X"A9",X"5A",X"95",X"5A",X"F5",
		X"AA",X"20",X"A2",X"FA",X"F7",X"B6",X"AA",X"AA",X"5B",X"6B",X"55",X"B5",X"AD",X"02",X"49",X"52",
		X"55",X"01",X"08",X"48",X"AA",X"52",X"D5",X"FD",X"77",X"55",X"AD",X"BB",X"DB",X"12",X"91",X"AA",
		X"AD",X"44",X"2A",X"49",X"55",X"22",X"AA",X"AA",X"AA",X"52",X"FF",X"FF",X"2A",X"25",X"AA",X"DA",
		X"6A",X"AD",X"2A",X"25",X"84",X"44",X"24",X"69",X"5B",X"AD",X"AA",X"DB",X"DB",X"AA",X"AA",X"52",
		X"6F",X"05",X"94",X"AA",X"AA",X"2A",X"49",X"AA",X"FA",X"5B",X"95",X"EA",X"ED",X"AE",X"AA",X"0A",
		X"B5",X"AA",X"04",X"52",X"B5",X"4A",X"22",X"48",X"DB",X"8A",X"54",X"A9",X"FF",X"AD",X"DB",X"DA",
		X"6E",X"15",X"48",X"A4",X"55",X"8A",X"D4",X"DA",X"ED",X"82",X"0A",X"92",X"52",X"52",X"25",X"B5",
		X"BD",X"E8",X"F6",X"56",X"5F",X"15",X"AA",X"AA",X"AA",X"57",X"68",X"15",X"12",X"95",X"54",X"55",
		X"D5",X"EA",X"77",X"B7",X"F6",X"55",X"AD",X"0A",X"51",X"15",X"AA",X"52",X"89",X"AA",X"88",X"D4",
		X"96",X"FE",X"95",X"EA",X"DE",X"EA",X"AD",X"54",X"55",X"44",X"92",X"4A",X"AB",X"54",X"12",X"49",
		X"54",X"A5",X"AA",X"F6",X"DB",X"96",X"EA",X"5B",X"5B",X"55",X"90",X"52",X"2B",X"89",X"5A",X"ED",
		X"AD",X"22",X"51",X"DB",X"5B",X"85",X"4A",X"2F",X"52",X"25",X"ED",X"45",X"5D",X"48",X"AA",X"CA",
		X"7F",X"A9",X"B6",X"A2",X"2B",X"80",X"B7",X"2A",X"7D",X"A0",X"96",X"D4",X"AA",X"4A",X"5F",X"BC",
		X"42",X"D4",X"AA",X"52",X"21",X"55",X"AD",X"DA",X"B5",X"6A",X"D5",X"7A",X"A9",X"A2",X"6F",X"4B",
		X"48",X"EA",X"6F",X"DB",X"12",X"54",X"4B",X"0A",X"41",X"DA",X"B6",X"AA",X"12",X"B5",X"57",X"55",
		X"A2",X"BE",X"05",X"BD",X"A2",X"EE",X"89",X"5E",X"91",X"BE",X"50",X"55",X"A9",X"1F",X"D4",X"55",
		X"D4",X"57",X"A8",X"04",X"D5",X"42",X"6A",X"AB",X"7E",X"95",X"56",X"41",X"6D",X"A0",X"6A",X"D5",
		X"6F",X"A5",X"16",X"55",X"2F",X"6A",X"EF",X"12",X"B7",X"04",X"52",X"29",X"55",X"A9",X"AA",X"D5",
		X"AD",X"42",X"55",X"B5",X"E2",X"D5",X"95",X"0D",X"12",X"B4",X"AA",X"DA",X"A5",X"BE",X"A5",X"82",
		X"88",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"4A",X"A5",X"4A",X"AD",X"56",X"AB",X"D5",
		X"AA",X"AA",X"FA",X"75",X"AB",X"02",X"10",X"A5",X"AA",X"55",X"F5",X"8A",X"22",X"D5",X"AD",X"AA",
		X"77",X"B7",X"EA",X"4A",X"00",X"AA",X"D5",X"6A",X"AD",X"13",X"29",X"55",X"2B",X"B5",X"5A",X"A5",
		X"F6",X"AF",X"5B",X"55",X"00",X"52",X"55",X"6B",X"57",X"29",X"52",X"95",X"AA",X"56",X"A7",X"5E",
		X"77",X"EF",X"5B",X"01",X"48",X"A5",X"DA",X"AF",X"94",X"8A",X"C4",X"6A",X"A5",X"56",X"AB",X"D6",
		X"EF",X"DE",X"05",X"80",X"8A",X"D4",X"5F",X"AA",X"0A",X"A4",X"AA",X"6A",X"9D",X"58",X"B7",X"FE",
		X"AD",X"15",X"80",X"14",X"FA",X"B5",X"5A",X"05",X"4A",X"95",X"5B",X"AB",X"5A",X"D5",X"FE",X"DB",
		X"05",X"A0",X"40",X"BD",X"FA",X"4A",X"15",X"A8",X"AA",X"F5",X"A2",X"55",X"AA",X"FB",X"DD",X"29",
		X"10",X"A0",X"D5",X"BE",X"B4",X"02",X"95",X"D4",X"A9",X"95",X"6A",X"E9",X"7B",X"BF",X"08",X"04",
		X"34",X"B9",X"2F",X"57",X"82",X"45",X"AD",X"F2",X"E1",X"62",X"F5",X"BE",X"5E",X"04",X"42",X"A6",
		X"B6",X"6B",X"95",X"12",X"A9",X"B2",X"5A",X"3D",X"5E",X"EB",X"D7",X"87",X"03",X"41",X"E5",X"EA",
		X"F1",X"A8",X"22",X"55",X"6A",X"9C",X"2E",X"57",X"AF",X"D7",X"E1",X"20",X"91",X"54",X"AB",X"AD",
		X"16",X"4A",X"B1",X"F0",X"78",X"BC",X"56",X"AF",X"4E",X"39",X"28",X"51",X"C3",X"93",X"1D",X"5A",
		X"54",X"A9",X"D1",X"E9",X"B4",X"3A",X"5D",X"AB",X"34",X"2A",X"2C",X"07",X"47",X"E5",X"70",X"5A",
		X"2C",X"16",X"57",X"7A",X"B5",X"5A",X"C7",X"86",X"E7",X"68",X"71",X"A8",X"51",X"C3",X"71",X"AC",
		X"1A",X"27",X"4E",X"17",X"1E",X"C7",X"87",X"63",X"9D",X"F1",X"58",X"72",X"8E",X"1C",X"E3",X"99",
		X"E1",X"38",X"9C",X"63",X"C7",X"31",X"8E",X"3A",X"E7",X"4C",X"63",X"1C",X"33",X"C6",X"E6",X"8C",
		X"63",X"CC",X"F2",X"54",X"78",X"1C",X"4E",X"1E",X"67",X"18",X"63",X"C6",X"B8",X"39",X"1B",X"87",
		X"63",X"E5",X"18",X"37",X"C6",X"F4",X"4C",X"8C",X"33",X"E3",X"38",X"E3",X"99",X"73",X"16",X"73",
		X"AC",X"33",X"C6",X"9D",X"E3",X"54",X"93",X"17",X"4E",X"E7",X"18",X"E3",X"E9",X"AC",X"D1",X"E1",
		X"58",X"E6",X"1C",X"1D",X"63",X"EA",X"58",X"39",X"C3",X"62",X"C6",X"B1",X"B1",X"52",X"8E",X"CD",
		X"84",X"71",X"E6",X"54",X"8E",X"8D",X"4A",X"96",X"59",X"19",X"E7",X"CC",X"19",X"C7",X"CA",X"71",
		X"72",X"66",X"CC",X"CC",X"CD",X"51",X"71",X"6E",X"9C",X"71",X"F1",X"70",X"72",X"63",X"AC",X"75",
		X"C6",X"99",X"38",X"76",X"A3",X"E2",X"C9",X"64",X"67",X"66",X"C6",X"CC",X"49",X"ED",X"98",X"61",
		X"6C",X"8C",X"16",X"E7",X"9C",X"31",X"66",X"8C",X"33",X"66",X"CE",X"64",X"E6",X"1C",X"39",X"CC",
		X"DC",X"38",X"67",X"86",X"67",X"CC",X"31",X"CE",X"31",X"26",X"8F",X"71",X"E6",X"C8",X"29",X"0F",
		X"33",X"66",X"CC",X"6E",X"AC",X"4C",X"1C",X"E6",X"66",X"29",X"63",X"9C",X"73",X"E6",X"9C",X"33",
		X"32",X"33",X"B3",X"1C",X"33",X"66",X"39",X"E6",X"8C",X"33",X"9C",X"71",X"CC",X"38",X"CF",X"8C",
		X"73",X"C6",X"38",X"67",X"C6",X"85",X"73",X"74",X"2C",X"C7",X"CE",X"18",X"AB",X"1A",X"B9",X"31",
		X"8D",X"53",X"CE",X"12",X"E7",X"38",X"E6",X"9C",X"4C",X"33",X"CD",X"38",X"CB",X"1C",X"63",X"9C",
		X"33",X"4B",X"6A",X"B3",X"C2",X"39",X"33",X"66",X"CE",X"94",X"69",X"4E",X"39",X"66",X"3C",X"33",
		X"47",X"76",X"27",X"2A",X"97",X"33",X"C5",X"1C",X"A7",X"32",X"39",X"66",X"56",X"C6",X"E6",X"A8",
		X"2A",X"3B",X"55",X"B2",X"31",X"9A",X"59",X"AE",X"96",X"C9",X"D0",X"AA",X"16",X"6B",X"D4",X"A8",
		X"55",X"A3",X"5A",X"95",X"AA",X"56",X"55",X"AA",X"AA",X"55",X"55",X"A5",X"AA",X"AA",X"AA",X"AA",
		X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"3A",X"9E",
		X"55",X"65",X"CC",X"A2",X"3A",X"CE",X"9C",X"19",X"5D",X"81",X"71",X"07",X"C7",X"CF",X"B8",X"3A",
		X"16",X"5D",X"E5",X"32",X"33",X"67",X"91",X"39",X"63",X"47",X"CE",X"98",X"D5",X"74",X"89",X"99",
		X"CB",X"32",X"C7",X"39",X"73",X"54",X"4A",X"33",X"63",X"9C",X"99",X"91",X"33",X"99",X"C5",X"73",
		X"62",X"2C",X"A6",X"67",X"DC",X"64",X"CE",X"C9",X"B2",X"99",X"CB",X"B1",X"31",X"8E",X"99",X"73",
		X"74",X"1C",X"57",X"E6",X"71",X"65",X"E6",X"A6",X"B9",X"AA",X"4A",X"3C",X"39",X"55",X"59",X"D3",
		X"81",X"9B",X"8B",X"63",X"EC",X"38",X"66",X"78",X"14",X"87",X"C3",X"71",X"74",X"1C",X"A6",X"E1",
		X"F0",X"E8",X"8C",X"1C",X"C7",X"CC",X"38",X"E6",X"AA",X"2A",X"C7",X"F1",X"78",X"1C",X"8F",X"E3",
		X"F1",X"68",X"BA",X"8A",X"C7",X"51",X"35",X"AD",X"AA",X"CE",X"F2",X"70",X"55",X"5D",X"8D",X"8B",
		X"A2",X"50",X"31",X"3A",X"CB",X"C5",X"A3",X"73",X"7D",X"BD",X"0E",X"03",X"A0",X"A2",X"1D",X"3F",
		X"AE",X"50",X"A1",X"E3",X"F5",X"7D",X"97",X"22",X"80",X"A8",X"EA",X"EE",X"56",X"15",X"05",X"95",
		X"FA",X"FC",X"BD",X"AE",X"1C",X"08",X"98",X"D4",X"A7",X"4F",X"17",X"8A",X"42",X"D5",X"EB",X"7B",
		X"D7",X"C5",X"40",X"20",X"9A",X"EE",X"AE",X"55",X"51",X"50",X"E2",X"DA",X"7D",X"FB",X"2E",X"0E",
		X"04",X"C4",X"AA",X"D7",X"AB",X"23",X"12",X"31",X"AD",X"DE",X"DD",X"B7",X"8B",X"02",X"82",X"E2",
		X"EA",X"5D",X"5D",X"0A",X"2A",X"38",X"F5",X"EA",X"5E",X"DF",X"E1",X"80",X"A0",X"54",X"BD",X"5E",
		X"5D",X"24",X"8A",X"54",X"AD",X"DE",X"DD",X"7D",X"C5",X"00",X"22",X"B8",X"BA",X"5B",X"17",X"15",
		X"51",X"54",X"B5",X"EB",X"BE",X"7E",X"15",X"05",X"88",X"68",X"75",X"BB",X"5A",X"85",X"0A",X"55",
		X"AA",X"6B",X"7F",X"FD",X"8A",X"0A",X"88",X"D0",X"6A",X"DD",X"55",X"55",X"14",X"A9",X"AA",X"EA",
		X"DD",X"DD",X"9D",X"0A",X"08",X"45",X"A9",X"D6",X"97",X"AB",X"54",X"8A",X"52",X"B5",X"FA",X"56",
		X"75",X"55",X"A2",X"2A",X"AA",X"54",X"55",X"55",X"55",X"D5",X"AA",X"AA",X"52",X"55",X"BD",X"AA",
		X"5B",X"B5",X"4A",X"15",X"AA",X"54",X"A5",X"4A",X"95",X"AA",X"55",X"AD",X"AA",X"52",X"55",X"55",
		X"AA",X"AA",X"AA",X"AA",X"55",X"55",X"45",X"95",X"AA",X"AA",X"6A",X"55",X"D5",X"AA",X"54",X"A9",
		X"5A",X"55",X"55",X"55",X"A9",X"52",X"B5",X"2A",X"55",X"AB",X"4A",X"55",X"95",X"AA",X"AA",X"56",
		X"55",X"55",X"55",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"55",X"A9",X"AA",X"AA",X"AA",X"CA",X"AA",
		X"54",X"A9",X"52",X"55",X"55",X"55",X"AB",X"54",X"A9",X"4A",X"55",X"AA",X"56",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"52",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"15",X"55",X"AB",X"56",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"38",X"3E",X"3C",X"7C",X"78",X"8E",X"73",X"F0",X"38",X"3C",X"0F",X"8F",X"C3",
		X"E1",X"6A",X"55",X"A9",X"72",X"91",X"6A",X"15",X"AB",X"4A",X"E5",X"70",X"74",X"87",X"F1",X"70",
		X"1C",X"C7",X"C3",X"83",X"87",X"C3",X"79",X"5C",X"1C",X"AB",X"AA",X"8B",X"C3",X"D5",X"1C",X"8B",
		X"63",X"D5",X"38",X"C5",X"A9",X"5A",X"B9",X"98",X"D5",X"E1",X"54",X"A5",X"E3",X"71",X"8A",X"C7",
		X"E1",X"38",X"AE",X"F2",X"70",X"5C",X"C3",X"63",X"8E",X"BA",X"2A",X"1E",X"1E",X"15",X"2D",X"9A",
		X"1A",X"AB",X"72",X"95",X"E3",X"75",X"AD",X"16",X"87",X"0A",X"19",X"3A",X"1E",X"8D",X"2A",X"D5",
		X"AA",X"7B",X"DD",X"5D",X"97",X"82",X"20",X"32",X"75",X"55",X"A5",X"A2",X"AA",X"AE",X"DE",X"7D",
		X"5F",X"C5",X"C0",X"20",X"56",X"8D",X"4B",X"95",X"4A",X"95",X"EA",X"76",X"BD",X"7F",X"C3",X"41",
		X"50",X"AA",X"56",X"55",X"A3",X"AA",X"54",X"55",X"F5",X"FA",X"FA",X"75",X"14",X"04",X"A6",X"56",
		X"B9",X"54",X"B1",X"4A",X"95",X"4A",X"D5",X"EB",X"7D",X"5D",X"0C",X"88",X"A2",X"4A",X"55",X"55",
		X"55",X"AA",X"AA",X"28",X"55",X"B5",X"FA",X"EE",X"55",X"15",X"0A",X"54",X"A4",X"6A",X"B5",X"6A",
		X"55",X"AA",X"54",X"AD",X"DE",X"F7",X"BB",X"8A",X"82",X"60",X"51",X"55",X"AD",X"AB",X"AA",X"16",
		X"55",X"55",X"F7",X"BA",X"BB",X"1A",X"15",X"81",X"A2",X"52",X"B5",X"5A",X"D5",X"2A",X"55",X"A9",
		X"56",X"AF",X"DF",X"55",X"A5",X"20",X"28",X"4A",X"55",X"AB",X"AA",X"6B",X"55",X"94",X"AA",X"DE",
		X"F5",X"DD",X"AA",X"02",X"44",X"91",X"AA",X"55",X"AB",X"55",X"A9",X"52",X"B5",X"6A",X"DD",X"EB",
		X"6A",X"0A",X"11",X"44",X"A5",X"AA",X"AA",X"5A",X"55",X"55",X"A5",X"AA",X"EA",X"5F",X"5D",X"55",
		X"8A",X"10",X"91",X"4A",X"55",X"EA",X"56",X"A9",X"52",X"A5",X"5A",X"BD",X"BE",X"5B",X"55",X"A1",
		X"A8",X"48",X"55",X"A5",X"AA",X"AA",X"55",X"95",X"AA",X"6A",X"55",X"BF",X"AA",X"2E",X"55",X"A1",
		X"2A",X"52",X"91",X"6A",X"95",X"AA",X"55",X"AB",X"54",X"AD",X"4A",X"95",X"EA",X"55",X"55",X"A9",
		X"AA",X"22",X"55",X"55",X"55",X"AD",X"AA",X"EA",X"5A",X"55",X"55",X"A9",X"AA",X"AA",X"55",X"95",
		X"2A",X"55",X"AA",X"56",X"A8",X"56",X"A5",X"6A",X"55",X"AA",X"54",X"AB",X"6A",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"A5",X"AA",X"AA",X"52",X"55",X"55",X"95",X"AA",X"6A",X"55",X"AD",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"CA",X"A3",X"F0",X"55",X"D1",X"AC",
		X"AA",X"1A",X"5F",X"05",X"73",X"1B",X"6A",X"71",X"71",X"AD",X"CC",X"43",X"B5",X"9C",X"4C",X"CB",
		X"74",X"D9",X"A8",X"5A",X"92",X"CA",X"4D",X"24",X"4E",X"AB",X"A5",X"74",X"8A",X"CC",X"62",X"A6",
		X"9D",X"56",X"5B",X"A5",X"46",X"6E",X"55",X"29",X"2D",X"BA",X"55",X"19",X"35",X"DB",X"B0",X"49",
		X"CE",X"AC",X"4C",X"B6",X"C9",X"A2",X"1A",X"4C",X"67",X"31",X"36",X"66",X"93",X"31",X"2F",X"8E",
		X"5E",X"71",X"3C",X"BA",X"C3",X"E5",X"3C",X"8E",X"E7",X"62",X"1C",X"8F",X"B3",X"2A",X"9E",X"59",
		X"31",X"CE",X"8E",X"D1",X"F1",X"A8",X"E2",X"C4",X"C5",X"0D",X"2B",X"87",X"1D",X"1D",X"8E",X"5A",
		X"39",X"EA",X"70",X"AA",X"D2",X"31",X"8E",X"1E",X"5D",X"3C",X"6A",X"74",X"74",X"8A",X"8B",X"79",
		X"74",X"AC",X"F2",X"38",X"D5",X"E1",X"B1",X"1A",X"0F",X"C7",X"39",X"3C",X"0E",X"D5",X"A8",X"AA",
		X"C5",X"A3",X"47",X"A7",X"2B",X"57",X"8F",X"8B",X"41",X"51",X"0E",X"8F",X"C7",X"2A",X"56",X"A5",
		X"7B",X"FD",X"ED",X"C1",X"81",X"88",X"C6",X"E5",X"95",X"8A",X"8A",X"54",X"BD",X"7A",X"BD",X"AF",
		X"0A",X"04",X"91",X"5A",X"DD",X"A9",X"18",X"2C",X"5A",X"D5",X"EB",X"F6",X"77",X"19",X"00",X"8A",
		X"EB",X"AE",X"45",X"05",X"47",X"47",X"AF",X"AE",X"EE",X"BF",X"70",X"40",X"B0",X"EA",X"D5",X"8A",
		X"43",X"A5",X"5A",X"55",X"AB",X"DD",X"FF",X"8A",X"80",X"90",X"CE",X"57",X"55",X"14",X"5A",X"EA",
		X"B8",X"54",X"DD",X"BF",X"2B",X"02",X"14",X"AA",X"77",X"55",X"28",X"71",X"AC",X"CA",X"A5",X"6B",
		X"DF",X"2F",X"22",X"20",X"AA",X"7D",X"D1",X"51",X"58",X"A9",X"AA",X"CA",X"D3",X"FD",X"BD",X"18",
		X"00",X"71",X"F9",X"54",X"A3",X"62",X"55",X"1A",X"97",X"EB",X"FA",X"7D",X"11",X"10",X"92",X"AE",
		X"4B",X"47",X"A5",X"AA",X"62",X"55",X"F5",X"FA",X"7B",X"15",X"02",X"42",X"75",X"AE",X"56",X"A5",
		X"4A",X"C5",X"AA",X"D6",X"F7",X"FB",X"A2",X"80",X"82",X"6A",X"55",X"5D",X"8B",X"AA",X"2A",X"AA",
		X"56",X"D7",X"F7",X"B5",X"A2",X"48",X"90",X"8A",X"52",X"BB",X"5A",X"95",X"AA",X"54",X"EF",X"FE",
		X"55",X"14",X"01",X"51",X"AA",X"AA",X"AE",X"AB",X"56",X"45",X"F5",X"BE",X"AB",X"22",X"42",X"50",
		X"A1",X"6A",X"B5",X"AA",X"55",X"AB",X"54",X"BF",X"AF",X"12",X"11",X"90",X"2A",X"6A",X"F5",X"6A",
		X"55",X"AD",X"52",X"7F",X"BF",X"8A",X"20",X"42",X"45",X"55",X"B5",X"AD",X"AA",X"AA",X"4A",X"F7",
		X"7D",X"8B",X"88",X"80",X"52",X"A9",X"6A",X"F5",X"AA",X"54",X"AD",X"DE",X"FD",X"AA",X"08",X"01",
		X"A5",X"AA",X"6A",X"DD",X"AA",X"55",X"A9",X"DE",X"FD",X"2A",X"0A",X"02",X"45",X"55",X"55",X"AF",
		X"AE",X"AA",X"4A",X"DD",X"77",X"2D",X"82",X"82",X"48",X"95",X"5A",X"DD",X"AA",X"55",X"A9",X"DE",
		X"BD",X"AA",X"40",X"41",X"A4",X"AA",X"D2",X"BD",X"5A",X"D5",X"AA",X"F7",X"BD",X"24",X"08",X"42",
		X"55",X"55",X"DD",X"E5",X"AA",X"2A",X"D5",X"F7",X"5D",X"06",X"82",X"A0",X"96",X"AA",X"57",X"AB",
		X"52",X"55",X"EA",X"7F",X"8F",X"82",X"10",X"54",X"A9",X"56",X"B7",X"4A",X"95",X"AA",X"F5",X"9F",
		X"E3",X"20",X"10",X"71",X"74",X"75",X"BA",X"AA",X"54",X"55",X"7F",X"3B",X"87",X"20",X"48",X"55",
		X"AD",X"56",X"97",X"4A",X"D5",X"FA",X"DD",X"E3",X"80",X"40",X"51",X"AD",X"CE",X"B5",X"2A",X"C6",
		X"AA",X"7F",X"9D",X"41",X"08",X"8A",X"55",X"75",X"9E",X"AA",X"52",X"D5",X"FB",X"3A",X"0E",X"42",
		X"84",X"4E",X"D5",X"BA",X"1C",X"8D",X"56",X"BF",X"6B",X"0E",X"02",X"21",X"A7",X"AE",X"7A",X"15",
		X"A5",X"AA",X"FF",X"79",X"0C",X"04",X"2A",X"1E",X"D7",X"5A",X"15",X"8E",X"F5",X"7E",X"1E",X"05",
		X"14",X"92",X"AE",X"5D",X"55",X"85",X"AA",X"DB",X"5F",X"0F",X"03",X"82",X"54",X"CF",X"D5",X"A5",
		X"48",X"D5",X"FB",X"D7",X"61",X"80",X"88",X"EA",X"75",X"71",X"89",X"A8",X"FA",X"FD",X"3C",X"04",
		X"28",X"38",X"7D",X"AE",X"16",X"28",X"56",X"BF",X"9F",X"07",X"01",X"61",X"AE",X"57",X"87",X"83",
		X"D2",X"F9",X"7B",X"35",X"04",X"04",X"AB",X"EF",X"5C",X"14",X"94",X"BA",X"FF",X"D5",X"50",X"40",
		X"A8",X"D7",X"AB",X"61",X"C1",X"E8",X"F7",X"8F",X"07",X"02",X"61",X"77",X"AF",X"8A",X"A0",X"D4",
		X"FD",X"3F",X"0E",X"00",X"C5",X"F5",X"75",X"99",X"88",X"D4",X"ED",X"7F",X"1C",X"00",X"A2",X"EB",
		X"EB",X"52",X"41",X"A9",X"BB",X"7F",X"1C",X"10",X"84",X"EB",X"CB",X"A5",X"48",X"B4",X"BE",X"3F",
		X"0E",X"04",X"C2",X"F6",X"B5",X"2A",X"28",X"B5",X"FE",X"1F",X"0D",X"10",X"E4",X"EA",X"B3",X"51",
		X"24",X"ED",X"FE",X"0F",X"0B",X"40",X"71",X"ED",X"5A",X"89",X"14",X"DF",X"FE",X"C3",X"01",X"84",
		X"BA",X"5E",X"55",X"A1",X"62",X"DF",X"FF",X"B0",X"00",X"11",X"AF",X"9E",X"2A",X"64",X"F1",X"BB",
		X"3F",X"1C",X"40",X"C1",X"A7",X"17",X"0D",X"AA",X"FC",X"ED",X"87",X"03",X"14",X"FC",X"78",X"15",
		X"0B",X"56",X"BF",X"FB",X"50",X"01",X"15",X"BD",X"BA",X"A2",X"42",X"ED",X"FD",X"17",X"0C",X"50",
		X"E2",X"57",X"AD",X"50",X"D4",X"DE",X"7F",X"B0",X"00",X"0B",X"7D",X"EA",X"42",X"25",X"FE",X"FC",
		X"83",X"06",X"68",X"D1",X"97",X"2D",X"A8",X"E2",X"5F",X"3F",X"B0",X"80",X"26",X"3F",X"D5",X"04",
		X"4E",X"FD",X"EE",X"83",X"04",X"B4",X"E8",X"97",X"2A",X"54",X"E9",X"77",X"57",X"04",X"A4",X"AA",
		X"BE",X"54",X"41",X"75",X"DF",X"5B",X"28",X"A0",X"4A",X"BD",X"2A",X"45",X"E9",X"D7",X"B7",X"82",
		X"40",X"B5",X"6A",X"95",X"8A",X"D2",X"AF",X"AF",X"05",X"41",X"74",X"DA",X"2A",X"2A",X"AA",X"DF",
		X"5D",X"05",X"8A",X"A8",X"56",X"57",X"A4",X"68",X"FD",X"EB",X"16",X"A0",X"48",X"DD",X"AA",X"05",
		X"AA",X"F6",X"D7",X"2D",X"A0",X"28",X"5B",X"55",X"15",X"B1",X"EA",X"AF",X"5B",X"40",X"54",X"D5",
		X"AA",X"2A",X"54",X"AD",X"7E",X"57",X"82",X"50",X"A5",X"5B",X"35",X"48",X"B5",X"EF",X"AE",X"44",
		X"44",X"55",X"AB",X"AA",X"82",X"5A",X"DF",X"5D",X"05",X"89",X"AA",X"BA",X"55",X"11",X"AA",X"DB",
		X"B7",X"2A",X"44",X"AA",X"5A",X"AD",X"42",X"D1",X"BA",X"77",X"55",X"90",X"A2",X"AA",X"AA",X"16",
		X"51",X"DD",X"B7",X"AB",X"A0",X"A8",X"54",X"55",X"95",X"2A",X"F5",X"EB",X"56",X"A1",X"0A",X"55",
		X"AB",X"54",X"AC",X"5E",X"DD",X"AA",X"A0",X"4A",X"5A",X"55",X"45",X"A9",X"EA",X"FA",X"5A",X"11",
		X"55",X"51",X"AD",X"A2",X"D4",X"AD",X"5B",X"D5",X"0A",X"15",X"A9",X"56",X"A9",X"6A",X"F5",X"AA",
		X"4B",X"55",X"11",X"A9",X"AA",X"AA",X"5A",X"55",X"D7",X"55",X"AA",X"0A",X"AA",X"4A",X"55",X"D5",
		X"AA",X"EA",X"55",X"AD",X"42",X"45",X"AA",X"54",X"AD",X"56",X"B5",X"6A",X"55",X"2A",X"54",X"A1",
		X"4A",X"D5",X"AA",X"5A",X"55",X"55",X"AD",X"88",X"2A",X"4A",X"55",X"55",X"DD",X"AA",X"AA",X"AA",
		X"52",X"51",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"4A",X"25",X"49",X"55",X"6D",X"55",X"55",
		X"55",X"55",X"B5",X"6E",X"EB",X"B7",X"52",X"55",X"55",X"D5",X"DB",X"56",X"AB",X"ED",X"EE",X"B6",
		X"AA",X"5A",X"DB",X"76",X"AD",X"25",X"A9",X"6A",X"AB",X"AA",X"AA",X"AA",X"2A",X"49",X"55",X"D5",
		X"5A",X"AB",X"22",X"25",X"55",X"55",X"4A",X"AA",X"B6",X"AA",X"AA",X"AA",X"AA",X"EF",X"AB",X"92",
		X"54",X"55",X"BB",X"AA",X"AA",X"AA",X"BE",X"55",X"A5",X"54",X"A9",X"AE",X"AA",X"5A",X"BD",X"52",
		X"29",X"49",X"24",X"89",X"24",X"AA",X"AA",X"24",X"0A",X"AA",X"54",X"08",X"52",X"AA",X"56",X"92",
		X"28",X"4A",X"55",X"24",X"22",X"29",X"85",X"A4",X"52",X"55",X"55",X"55",X"95",X"BA",X"5F",X"D5",
		X"F6",X"F7",X"DD",X"B6",X"AA",X"6E",X"D5",X"6E",X"6B",X"55",X"B5",X"BA",X"5D",X"25",X"92",X"54",
		X"7F",X"B7",X"0A",X"AA",X"DA",X"5B",X"15",X"59",X"EF",X"B7",X"B6",X"4A",X"95",X"BA",X"55",X"25",
		X"54",X"AD",X"DF",X"AA",X"8A",X"48",X"55",X"95",X"28",X"59",X"AB",X"56",X"BD",X"AD",X"55",X"15",
		X"55",X"22",X"09",X"20",X"49",X"25",X"85",X"90",X"44",X"52",X"B5",X"94",X"14",X"8A",X"44",X"AA",
		X"52",X"88",X"10",X"A5",X"DA",X"BD",X"EB",X"DE",X"7B",X"B7",X"6B",X"BB",X"BD",X"6B",X"AB",X"EA",
		X"76",X"55",X"55",X"54",X"B7",X"55",X"50",X"7D",X"FF",X"B6",X"B6",X"FB",X"BD",X"B5",X"D4",X"6D",
		X"AB",X"90",X"52",X"55",X"10",X"00",X"94",X"94",X"12",X"88",X"2A",X"95",X"A4",X"54",X"6B",X"DB",
		X"AA",X"6A",X"FB",X"77",X"BB",X"FD",X"2B",X"00",X"00",X"00",X"00",X"00",X"49",X"B5",X"AA",X"94",
		X"52",X"55",X"55",X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"EF",X"15",X"02",X"00",X"82",X"10",
		X"52",X"DD",X"BF",X"5B",X"95",X"24",X"11",X"21",X"69",X"FB",X"FF",X"FD",X"FF",X"FF",X"7D",X"6F",
		X"25",X"00",X"00",X"00",X"00",X"00",X"B2",X"DB",X"B5",X"55",X"09",X"00",X"00",X"D2",X"76",X"BF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"0B",X"00",X"00",X"00",X"00",X"50",X"FB",X"7F",X"B7",X"55",X"09",
		X"00",X"00",X"D4",X"BD",X"F7",X"FF",X"FF",X"FF",X"FF",X"5F",X"00",X"00",X"00",X"00",X"00",X"B4",
		X"FF",X"DE",X"96",X"04",X"00",X"00",X"80",X"BA",X"F7",X"FF",X"FF",X"FF",X"FF",X"97",X"00",X"00",
		X"00",X"00",X"00",X"BA",X"FF",X"BD",X"AD",X"02",X"00",X"00",X"20",X"7B",X"DF",X"FF",X"FF",X"FF",
		X"FF",X"0B",X"00",X"00",X"00",X"00",X"40",X"FB",X"7F",X"DF",X"55",X"01",X"00",X"00",X"90",X"7B",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"05",X"00",X"00",X"00",X"00",X"D0",X"FF",X"FB",X"DD",X"96",X"00",
		X"00",X"00",X"D4",X"BB",X"FF",X"FF",X"FF",X"FF",X"5F",X"00",X"00",X"00",X"00",X"00",X"BA",X"FF",
		X"DF",X"DB",X"4A",X"00",X"00",X"00",X"79",X"EF",X"FF",X"FF",X"FF",X"FF",X"17",X"00",X"00",X"00",
		X"00",X"80",X"F6",X"FF",X"F7",X"B6",X"09",X"00",X"00",X"80",X"BA",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"4B",X"00",X"00",X"00",X"00",X"80",X"EE",X"FF",X"F7",X"6D",X"05",X"00",X"00",X"80",X"BA",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"17",X"01",X"00",X"00",X"00",X"80",X"FA",X"BF",X"FF",X"B6",X"25",X"00",
		X"00",X"00",X"EA",X"BB",X"FF",X"FF",X"FF",X"FF",X"BF",X"08",X"00",X"00",X"00",X"00",X"E8",X"FE",
		X"7F",X"AF",X"2B",X"01",X"00",X"00",X"A0",X"FD",X"DE",X"FF",X"FF",X"FF",X"FF",X"2B",X"00",X"00",
		X"00",X"00",X"80",X"EE",X"FF",X"BE",X"6D",X"49",X"00",X"00",X"00",X"74",X"BF",X"F7",X"FF",X"FF",
		X"FF",X"7F",X"05",X"00",X"00",X"00",X"00",X"A0",X"FD",X"7E",X"6F",X"AB",X"12",X"00",X"00",X"00",
		X"FA",X"7D",X"EF",X"FF",X"FF",X"FF",X"7F",X"05",X"00",X"00",X"00",X"00",X"50",X"FB",X"7E",X"77",
		X"AD",X"12",X"02",X"00",X"00",X"F4",X"7B",X"F7",X"FF",X"FF",X"FF",X"FF",X"0D",X"00",X"00",X"00",
		X"00",X"40",X"ED",X"FD",X"DE",X"AE",X"2A",X"01",X"00",X"00",X"C8",X"DF",X"BB",X"FF",X"FF",X"FF",
		X"FF",X"DF",X"00",X"00",X"00",X"00",X"00",X"54",X"DF",X"EF",X"ED",X"6A",X"29",X"00",X"00",X"00",
		X"F5",X"7B",X"F7",X"FF",X"FF",X"FF",X"FF",X"6F",X"00",X"00",X"00",X"00",X"00",X"EA",X"EE",X"EF",
		X"6E",X"AB",X"4A",X"00",X"00",X"80",X"EC",X"DF",X"DD",X"FF",X"FF",X"FF",X"FF",X"DF",X"00",X"00",
		X"00",X"00",X"00",X"64",X"EF",X"F7",X"ED",X"D6",X"2A",X"01",X"00",X"00",X"B2",X"7F",X"B7",X"EF",
		X"FF",X"FF",X"FF",X"FF",X"0B",X"00",X"00",X"00",X"00",X"90",X"FA",X"7E",X"DF",X"AE",X"AD",X"12",
		X"00",X"00",X"A0",X"F6",X"BB",X"BD",X"FF",X"FF",X"FF",X"FF",X"DF",X"00",X"00",X"00",X"00",X"00",
		X"52",X"EF",X"F7",X"BB",X"AD",X"55",X"22",X"00",X"00",X"68",X"BF",X"DB",X"FB",X"FF",X"FF",X"FF",
		X"FF",X"5B",X"00",X"00",X"00",X"00",X"80",X"74",X"EF",X"BF",X"DB",X"56",X"55",X"02",X"00",X"00",
		X"D6",X"F7",X"76",X"FF",X"FF",X"FF",X"FF",X"FF",X"0D",X"00",X"00",X"00",X"00",X"40",X"BA",X"BF",
		X"DF",X"6D",X"AD",X"25",X"21",X"00",X"00",X"6A",X"DF",X"ED",X"FB",X"FF",X"FF",X"FF",X"FF",X"2D",
		X"00",X"00",X"00",X"00",X"80",X"F4",X"FD",X"7B",X"DB",X"5A",X"4B",X"41",X"00",X"00",X"D4",X"BE",
		X"BB",X"EF",X"FF",X"FF",X"FF",X"FF",X"37",X"01",X"00",X"00",X"00",X"00",X"D2",X"F7",X"F7",X"B6",
		X"AD",X"55",X"09",X"00",X"00",X"C8",X"F6",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"DF",X"00",X"00",
		X"00",X"00",X"00",X"D2",X"FB",X"BB",X"6D",X"DB",X"AA",X"04",X"00",X"00",X"AA",X"6E",X"EF",X"FD",
		X"FF",X"FF",X"FF",X"FF",X"2B",X"00",X"00",X"00",X"00",X"90",X"BE",X"DF",X"6E",X"DB",X"B5",X"04",
		X"01",X"00",X"A4",X"6A",X"F7",X"FE",X"FD",X"FF",X"FF",X"FF",X"DF",X"00",X"00",X"00",X"00",X"00",
		X"D9",X"FB",X"B6",X"DD",X"6E",X"25",X"01",X"04",X"40",X"54",X"ED",X"DE",X"EF",X"FF",X"FF",X"FF",
		X"FF",X"1B",X"00",X"00",X"00",X"01",X"20",X"DD",X"BD",X"ED",X"EE",X"B6",X"14",X"44",X"00",X"10",
		X"2A",X"7B",X"EF",X"FD",X"FF",X"FF",X"FF",X"FF",X"2D",X"00",X"00",X"00",X"00",X"20",X"DD",X"BD",
		X"ED",X"76",X"57",X"25",X"44",X"80",X"00",X"4A",X"DD",X"BD",X"F7",X"FF",X"FF",X"FF",X"FF",X"5B",
		X"00",X"00",X"00",X"00",X"40",X"DA",X"BD",X"DB",X"DD",X"6D",X"95",X"10",X"81",X"00",X"44",X"D9",
		X"DD",X"BB",X"FF",X"FF",X"FF",X"FF",X"BF",X"05",X"00",X"00",X"00",X"00",X"C8",X"F6",X"EE",X"EE",
		X"EE",X"5A",X"09",X"11",X"02",X"80",X"50",X"DD",X"BD",X"FB",X"FF",X"FF",X"FF",X"FF",X"B7",X"04",
		X"00",X"00",X"00",X"00",X"B2",X"7D",X"77",X"BB",X"BB",X"55",X"42",X"08",X"81",X"00",X"94",X"DD",
		X"77",X"F7",X"FF",X"FF",X"DF",X"FF",X"B7",X"02",X"00",X"00",X"00",X"00",X"D2",X"DE",X"BB",X"DD",
		X"DD",X"9A",X"04",X"21",X"42",X"00",X"A2",X"DA",X"7B",X"BB",X"FF",X"FF",X"FF",X"FB",X"BF",X"0D",
		X"00",X"00",X"00",X"00",X"88",X"B6",X"EF",X"EE",X"76",X"5B",X"93",X"10",X"24",X"82",X"00",X"A9",
		X"EE",X"BB",X"BB",X"FF",X"FF",X"FF",X"FB",X"6F",X"05",X"00",X"00",X"00",X"00",X"A4",X"F6",X"DE",
		X"6E",X"BB",X"6D",X"49",X"08",X"22",X"81",X"80",X"54",X"7D",X"EF",X"EE",X"FF",X"FF",X"7F",X"FF",
		X"BD",X"0A",X"00",X"00",X"80",X"40",X"50",X"B5",X"77",X"B7",X"ED",X"B6",X"2A",X"21",X"10",X"89",
		X"08",X"22",X"B5",X"F7",X"DD",X"DE",X"FF",X"FF",X"DF",X"FF",X"B6",X"04",X"00",X"00",X"00",X"81",
		X"A8",X"FA",X"EE",X"B6",X"ED",X"B6",X"12",X"81",X"90",X"54",X"08",X"A1",X"DA",X"7E",X"DB",X"F6",
		X"FF",X"FF",X"7F",X"FF",X"B7",X"02",X"00",X"00",X"80",X"00",X"A1",X"F6",X"EE",X"B6",X"6D",X"BB",
		X"4A",X"02",X"21",X"A9",X"84",X"08",X"D5",X"EE",X"6D",X"BB",X"FF",X"FF",X"FF",X"DF",X"7F",X"8D",
		X"00",X"00",X"00",X"10",X"08",X"D5",X"DE",X"DB",X"B6",X"6D",X"AB",X"22",X"08",X"89",X"4A",X"42",
		X"48",X"6A",X"77",X"6F",X"F7",X"FF",X"FF",X"FF",X"FD",X"BB",X"12",X"00",X"00",X"00",X"08",X"44",
		X"B5",X"FB",X"6E",X"5B",X"6B",X"55",X"09",X"82",X"48",X"2A",X"89",X"24",X"B5",X"FB",X"EE",X"DE",
		X"FF",X"FF",X"FF",X"EF",X"B7",X"0A",X"00",X"00",X"00",X"04",X"92",X"AA",X"BB",X"77",X"5B",X"6B",
		X"55",X"85",X"08",X"22",X"49",X"25",X"89",X"54",X"ED",X"BE",X"F7",X"FE",X"FF",X"FF",X"BF",X"6F",
		X"95",X"00",X"00",X"00",X"80",X"88",X"54",X"BB",X"F7",X"EE",X"56",X"AB",X"4A",X"22",X"82",X"48",
		X"2A",X"95",X"92",X"52",X"DB",X"EF",X"7D",X"FF",X"FF",X"DF",X"BF",X"5B",X"25",X"00",X"00",X"00",
		X"20",X"92",X"AA",X"ED",X"BB",X"77",X"AB",X"96",X"12",X"11",X"41",X"44",X"2A",X"95",X"24",X"A9",
		X"EA",X"BE",X"77",X"F7",X"EF",X"FF",X"BF",X"6F",X"95",X"00",X"00",X"20",X"44",X"52",X"B5",X"7D",
		X"DF",X"77",X"AD",X"AA",X"24",X"42",X"20",X"44",X"94",X"94",X"24",X"24",X"55",X"6D",X"77",X"BB",
		X"F7",X"FF",X"FB",X"EF",X"AD",X"42",X"00",X"20",X"44",X"92",X"B2",X"DA",X"7B",X"77",X"AB",X"2A",
		X"89",X"08",X"10",X"10",X"92",X"54",X"29",X"11",X"91",X"D4",X"F6",X"B6",X"BD",X"FF",X"FF",X"FF",
		X"BF",X"6F",X"55",X"02",X"41",X"48",X"92",X"AA",X"6A",X"BB",X"5B",X"AB",X"2A",X"84",X"00",X"81",
		X"10",X"91",X"24",X"49",X"24",X"12",X"55",X"B5",X"DD",X"FD",X"FE",X"FB",X"FF",X"FF",X"EF",X"56",
		X"12",X"08",X"08",X"91",X"A4",X"AA",X"AA",X"5A",X"55",X"95",X"44",X"84",X"20",X"22",X"25",X"91",
		X"A4",X"24",X"89",X"90",X"AA",X"DB",X"F7",X"FE",X"EF",X"BF",X"FF",X"FF",X"BB",X"55",X"44",X"40",
		X"88",X"24",X"49",X"55",X"55",X"AD",X"AA",X"24",X"22",X"88",X"10",X"11",X"91",X"28",X"55",X"8A",
		X"20",X"A8",X"DA",X"BD",X"DD",X"FB",X"FF",X"FD",X"EF",X"FF",X"6F",X"15",X"01",X"21",X"44",X"22",
		X"A9",X"B6",X"5D",X"AB",X"AA",X"24",X"12",X"11",X"49",X"55",X"55",X"55",X"55",X"41",X"00",X"D2",
		X"F6",X"B6",X"FD",X"FF",X"BD",X"DF",X"FF",X"DF",X"2A",X"80",X"00",X"21",X"08",X"A9",X"EE",X"5B",
		X"55",X"52",X"89",X"00",X"00",X"49",X"A5",X"A4",X"6A",X"5B",X"01",X"00",X"54",X"F7",X"ED",X"FE",
		X"FF",X"7F",X"EF",X"FF",X"7F",X"21",X"90",X"04",X"02",X"B4",X"7E",X"AF",X"EB",X"5E",X"05",X"80",
		X"10",X"09",X"50",X"F5",X"56",X"55",X"55",X"00",X"00",X"68",X"B7",X"FD",X"FF",X"DF",X"DD",X"FF",
		X"BD",X"2B",X"10",X"00",X"00",X"20",X"AE",X"DB",X"DB",X"57",X"85",X"50",X"10",X"92",X"6D",X"5F",
		X"DF",X"DB",X"14",X"02",X"00",X"B0",X"B6",X"FF",X"BF",X"BB",X"7D",X"EF",X"FF",X"FF",X"05",X"00",
		X"00",X"00",X"E2",X"31",X"FF",X"AE",X"30",X"01",X"04",X"34",X"D9",X"EB",X"6F",X"57",X"25",X"20",
		X"40",X"D0",X"5E",X"FF",X"FD",X"D6",X"DD",X"7B",X"FF",X"FF",X"FF",X"40",X"00",X"00",X"20",X"BC",
		X"FE",X"A7",X"16",X"04",X"00",X"28",X"CB",X"7F",X"BD",X"53",X"01",X"02",X"21",X"5A",X"F3",X"7A",
		X"AB",X"B5",X"AE",X"F7",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"93",X"FF",X"7F",X"58",X"40",
		X"00",X"84",X"B6",X"FF",X"7D",X"55",X"02",X"40",X"A4",X"BA",X"EB",X"69",X"85",X"4A",X"5E",X"FF",
		X"FE",X"FF",X"FF",X"BF",X"0F",X"00",X"00",X"80",X"95",X"7F",X"3F",X"2C",X"00",X"00",X"51",X"AF",
		X"7F",X"BD",X"A4",X"00",X"84",X"54",X"B7",X"BB",X"5A",X"20",X"A2",X"F5",X"F7",X"BF",X"FF",X"EF",
		X"DF",X"AB",X"01",X"00",X"00",X"AC",X"FA",X"FB",X"A1",X"00",X"00",X"0A",X"7B",X"FD",X"FA",X"28",
		X"81",X"80",X"8A",X"AE",X"BE",X"5A",X"94",X"A8",X"EA",X"FB",X"F7",X"BF",X"FF",X"EF",X"2F",X"07",
		X"00",X"00",X"30",X"FB",X"F9",X"C3",X"01",X"00",X"14",X"D6",X"7E",X"FD",X"B4",X"40",X"81",X"88",
		X"56",X"AF",X"AE",X"94",X"58",X"75",X"FB",X"FB",X"FB",X"BF",X"FF",X"BE",X"4D",X"00",X"00",X"80",
		X"F8",X"EB",X"AB",X"06",X"00",X"04",X"34",X"FD",X"F6",X"BA",X"42",X"20",X"41",X"A5",X"D7",X"AD",
		X"0A",X"85",X"5A",X"FB",X"FE",X"7E",X"F7",X"FD",X"EF",X"6F",X"0B",X"00",X"00",X"C0",X"F8",X"77",
		X"59",X"06",X"00",X"90",X"A9",X"DE",X"6F",X"95",X"22",X"08",X"54",X"5D",X"5D",X"6B",X"41",X"A0",
		X"69",X"EF",X"BF",X"DB",X"ED",X"ED",X"F7",X"FF",X"75",X"02",X"00",X"00",X"0C",X"FF",X"8F",X"42",
		X"08",X"00",X"69",X"BD",X"7B",X"5D",X"09",X"08",X"49",X"D5",X"EE",X"55",X"85",X"20",X"52",X"BB",
		X"FF",X"DD",X"AE",X"ED",X"DD",X"FF",X"FF",X"DA",X"00",X"00",X"00",X"C3",X"FB",X"A7",X"01",X"08",
		X"02",X"A9",X"EF",X"57",X"4D",X"22",X"08",X"52",X"BB",X"DB",X"5A",X"12",X"40",X"B4",X"7D",X"77",
		X"77",X"AB",X"B6",X"EF",X"FF",X"FB",X"AF",X"2A",X"00",X"00",X"70",X"3C",X"FF",X"38",X"00",X"20",
		X"34",X"F5",X"7E",X"AD",X"90",X"10",X"91",X"D4",X"BE",X"5B",X"29",X"08",X"51",X"DA",X"F7",X"B6",
		X"B6",X"76",X"ED",X"FE",X"FD",X"7B",X"AB",X"34",X"00",X"00",X"68",X"3C",X"6E",X"35",X"00",X"50",
		X"54",X"D5",X"DA",X"AD",X"22",X"44",X"52",X"A9",X"EA",X"6E",X"4B",X"10",X"92",X"AA",X"F5",X"DE",
		X"5D",X"DB",X"EE",X"DE",X"FB",X"FF",X"55",X"A9",X"0A",X"00",X"00",X"8F",X"E3",X"5A",X"87",X"00",
		X"44",X"55",X"55",X"DD",X"AD",X"08",X"49",X"8A",X"A4",X"BA",X"DB",X"AA",X"02",X"A1",X"AA",X"B5",
		X"DE",X"DE",X"B6",X"BB",X"F7",X"EE",X"EF",X"96",X"4A",X"2D",X"00",X"00",X"69",X"38",X"DA",X"6A",
		X"10",X"A2",X"94",X"48",X"B5",X"AD",X"92",X"94",X"92",X"48",X"DA",X"B6",X"D5",X"B6",X"00",X"D4",
		X"EA",X"D4",X"FB",X"6D",X"B5",X"BB",X"EB",X"7E",X"EF",X"AA",X"52",X"05",X"00",X"A0",X"A4",X"50",
		X"D5",X"8A",X"44",X"95",X"44",X"52",X"55",X"25",X"55",X"55",X"A9",X"AA",X"AA",X"52",X"55",X"2B",
		X"54",X"DB",X"55",X"BA",X"56",X"D5",X"E2",X"E7",X"AF",X"5F",X"7D",X"DD",X"6A",X"55",X"55",X"40",
		X"20",X"84",X"A0",X"54",X"95",X"52",X"55",X"52",X"AA",X"4A",X"A9",X"AA",X"52",X"2A",X"A5",X"54",
		X"55",X"55",X"55",X"A5",X"AA",X"AA",X"D6",X"AA",X"AA",X"DE",X"BA",X"BD",X"ED",X"EE",X"B6",X"B6",
		X"D6",X"AA",X"2A",X"11",X"10",X"42",X"10",X"29",X"89",X"52",X"2A",X"A9",X"AA",X"AA",X"D5",X"AA",
		X"4A",X"55",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"B5",X"FA",X"56",X"6B",X"15",X"95",X"4A",X"A9",
		X"6A",X"AD",X"56",X"55",X"55",X"55",X"6F",X"5B",X"AB",X"24",X"49",X"42",X"44",X"08",X"11",X"22",
		X"24",X"91",X"A4",X"52",X"95",X"6A",X"B5",X"D6",X"AD",X"DA",X"5A",X"55",X"A9",X"92",X"4A",X"55",
		X"D5",X"F6",X"7B",X"77",X"BB",X"AD",X"B5",X"B5",X"B6",X"56",X"55",X"4A",X"AA",X"54",X"A9",X"AA",
		X"12",X"42",X"04",X"21",X"11",X"A5",X"54",X"AA",X"AA",X"AA",X"AA",X"D6",X"6D",X"B5",X"56",X"55",
		X"95",X"AA",X"AA",X"AA",X"6A",X"BD",X"AD",X"6D",X"AB",X"2D",X"A5",X"94",X"52",X"A9",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"4A",X"91",X"A4",X"A4",X"54",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"B5",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"C7",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"55",
		X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"6A",X"69",X"55",X"95",X"AA",X"AA",X"AA",X"2A",X"9A",X"96",X"AA",X"74",X"69",X"D1",X"B4",
		X"2A",X"AB",X"2A",X"B5",X"E8",X"AA",X"3C",X"5C",X"AC",X"54",X"D3",X"D2",X"D2",X"D1",X"D2",X"AA",
		X"5A",X"5C",X"2C",X"55",X"55",X"AD",X"52",X"55",X"55",X"A9",X"AA",X"AA",X"D2",X"07",X"0F",X"87",
		X"C3",X"C3",X"A9",X"CA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"9D",X"AA",X"AA",X"EA",X"B0",X"AA",
		X"74",X"AA",X"5A",X"AA",X"56",X"1D",X"4B",X"E3",X"E1",X"E1",X"45",X"E3",X"E1",X"E1",X"C5",X"51",
		X"1D",X"9E",X"D1",X"E1",X"E1",X"71",X"3C",X"A6",X"1C",X"9D",X"78",X"78",X"78",X"3C",X"9C",X"4A",
		X"4D",X"79",X"71",X"8E",X"A9",X"C0",X"C7",X"CA",X"E3",X"E1",X"E1",X"91",X"0F",X"3E",X"6C",X"39",
		X"1C",X"0F",X"8F",X"C3",X"C3",X"59",X"1C",X"8F",X"E3",X"F0",X"68",X"78",X"78",X"78",X"78",X"38",
		X"36",X"56",X"A5",X"87",X"47",X"4E",X"55",X"8D",X"75",X"38",X"1E",X"1E",X"5E",X"A8",X"C7",X"E1",
		X"38",X"2E",X"3C",X"0E",X"CF",X"70",X"0E",X"E7",X"38",X"1E",X"3E",X"1C",X"CF",X"E8",X"E2",X"E2",
		X"CC",X"1C",X"17",X"1E",X"1F",X"7C",X"C8",X"C3",X"43",X"7B",X"78",X"3C",X"1C",X"1E",X"C7",X"31",
		X"87",X"87",X"87",X"C3",X"87",X"6D",X"38",X"4E",X"3C",X"EA",X"C1",X"E3",X"F0",X"F0",X"C3",X"63",
		X"1C",X"1E",X"FC",X"E0",X"C1",X"87",X"0F",X"C7",X"C1",X"87",X"43",X"0F",X"F3",X"F0",X"C1",X"71",
		X"1C",X"87",X"CB",X"78",X"78",X"38",X"1E",X"3E",X"3C",X"1C",X"77",X"E0",X"E1",X"83",X"0F",X"3E",
		X"7C",X"C2",X"87",X"3E",X"AC",X"71",X"F8",X"E0",X"C3",X"71",X"0E",X"9E",X"C3",X"63",X"4E",X"F2",
		X"0A",X"8F",X"C3",X"31",X"3C",X"8E",X"74",X"E0",X"C3",X"C3",X"F0",X"78",X"78",X"0C",X"0F",X"0F",
		X"AF",X"F0",X"D8",X"0B",X"CF",X"E1",X"C1",X"47",X"0F",X"2F",X"1E",X"1E",X"5E",X"F0",X"C2",X"87",
		X"F0",X"C1",X"0F",X"78",X"54",X"A5",X"83",X"AB",X"78",X"A8",X"0F",X"1E",X"7C",X"F8",X"E0",X"63",
		X"87",X"57",X"FC",X"F0",X"D1",X"96",X"8B",X"2D",X"79",X"A8",X"8B",X"6A",X"68",X"54",X"95",X"0A",
		X"4B",X"85",X"1C",X"38",X"0C",X"EA",X"E0",X"E1",X"AA",X"E3",X"97",X"BF",X"FA",X"E9",X"D3",X"D2",
		X"A9",X"A5",X"0B",X"1F",X"3E",X"F4",X"AA",X"D3",X"BA",X"5A",X"DB",X"FA",X"F2",X"BA",X"72",X"71",
		X"41",X"83",X"42",X"21",X"50",X"A0",X"40",X"41",X"42",X"41",X"52",X"D1",X"B4",X"CE",X"AD",X"AE",
		X"74",X"30",X"21",X"54",X"C4",X"55",X"F4",X"F0",X"43",X"8F",X"0F",X"AF",X"FA",X"AA",X"16",X"9A",
		X"AA",X"BB",X"7C",X"A9",X"72",X"F8",X"C5",X"2F",X"7E",X"F4",X"FB",X"F1",X"A7",X"2F",X"BF",X"7A",
		X"BB",X"17",X"79",X"E1",X"85",X"05",X"02",X"0A",X"B6",X"A8",X"00",X"22",X"55",X"A5",X"40",X"45",
		X"D7",X"1E",X"7A",X"F0",X"0F",X"FE",X"F0",X"C3",X"0F",X"0F",X"2F",X"74",X"C0",X"05",X"DB",X"A2",
		X"85",X"2E",X"B4",X"AA",X"EA",X"AD",X"6F",X"ED",X"DA",X"6E",X"FB",X"CB",X"1F",X"BD",X"D6",X"3F",
		X"F8",X"81",X"07",X"40",X"00",X"05",X"A9",X"00",X"06",X"58",X"A1",X"8A",X"14",X"91",X"5A",X"EA",
		X"D2",X"4B",X"B7",X"BD",X"6E",X"7B",X"FD",X"BF",X"FF",X"E1",X"0F",X"18",X"80",X"5B",X"FC",X"01",
		X"0A",X"F8",X"AA",X"2E",X"68",X"41",X"5F",X"ED",X"2A",X"55",X"AA",X"BD",X"ED",X"7B",X"F7",X"DE",
		X"F6",X"FE",X"BF",X"FF",X"3F",X"C0",X"01",X"7F",X"C9",X"07",X"40",X"C0",X"FF",X"11",X"00",X"F8",
		X"ED",X"1F",X"00",X"3C",X"F8",X"A7",X"13",X"D2",X"5F",X"FE",X"D0",X"AF",X"F6",X"CB",X"FF",X"0F",
		X"70",X"80",X"7F",X"C0",X"03",X"F0",X"E1",X"3F",X"00",X"02",X"FE",X"4B",X"0B",X"80",X"AF",X"F6",
		X"02",X"48",X"F4",X"AF",X"54",X"52",X"7F",X"EB",X"56",X"DF",X"FA",X"1F",X"80",X"03",X"FE",X"03",
		X"08",X"C0",X"3F",X"3D",X"00",X"F8",X"F9",X"0F",X"00",X"A5",X"FF",X"41",X"11",X"C0",X"4F",X"3F",
		X"A0",X"7E",X"F5",X"85",X"DD",X"DF",X"6E",X"FD",X"01",X"E0",X"C1",X"7F",X"00",X"0C",X"F8",X"0F",
		X"A8",X"80",X"FF",X"50",X"05",X"E8",X"5F",X"AA",X"00",X"BD",X"F8",X"03",X"AC",X"F6",X"3D",X"E0",
		X"D7",X"BF",X"AA",X"BB",X"FE",X"03",X"E0",X"81",X"FF",X"00",X"1C",X"F8",X"0F",X"80",X"93",X"FE",
		X"03",X"B0",X"E2",X"BF",X"80",X"0A",X"DB",X"2D",X"40",X"FA",X"ED",X"15",X"AA",X"FF",X"6E",X"AD",
		X"ED",X"FF",X"03",X"C0",X"87",X"FF",X"02",X"E0",X"D2",X"3F",X"00",X"F8",X"AA",X"2F",X"00",X"DE",
		X"DA",X"0E",X"80",X"BB",X"E0",X"03",X"AE",X"2F",X"5D",X"69",X"FF",X"95",X"7E",X"6D",X"FF",X"07",
		X"80",X"1F",X"FA",X"07",X"80",X"BF",X"F0",X"03",X"C0",X"7F",X"E4",X"02",X"E0",X"7F",X"91",X"44",
		X"B0",X"7E",X"41",X"8B",X"76",X"3F",X"A9",X"6E",X"DF",X"57",X"DB",X"FE",X"7F",X"00",X"F8",X"07",
		X"FE",X"00",X"E0",X"1F",X"5A",X"00",X"E0",X"FF",X"02",X"29",X"50",X"FF",X"03",X"A8",X"92",X"BA",
		X"2D",X"D4",X"DE",X"5A",X"5B",X"F5",X"EF",X"DE",X"BA",X"FF",X"03",X"00",X"FE",X"E0",X"07",X"00",
		X"F8",X"5F",X"90",X"05",X"A0",X"FF",X"8A",X"24",X"25",X"D4",X"BB",X"40",X"2A",X"55",X"ED",X"55",
		X"AD",X"AD",X"76",X"B7",X"FE",X"6D",X"FD",X"FF",X"00",X"00",X"FE",X"21",X"D3",X"00",X"80",X"FF",
		X"15",X"4A",X"01",X"64",X"FF",X"16",X"91",X"88",X"A8",X"7B",X"15",X"91",X"AA",X"BE",X"5B",X"55",
		X"D5",X"EE",X"B7",X"DA",X"6D",X"F7",X"0F",X"00",X"C0",X"37",X"5A",X"0B",X"00",X"A0",X"FF",X"2A",
		X"89",X"22",X"A2",X"76",X"B7",X"42",X"A4",X"2A",X"48",X"ED",X"2B",X"AA",X"D5",X"5A",X"6B",X"7B",
		X"5B",X"B7",X"DB",X"EE",X"FB",X"0B",X"00",X"80",X"5D",X"2A",X"55",X"01",X"00",X"DB",X"AB",X"54",
		X"A6",X"22",X"54",X"6D",X"A5",X"AA",X"2A",X"01",X"D8",X"7D",X"55",X"AB",X"4A",X"ED",X"ED",X"6D",
		X"DB",X"B6",X"F7",X"76",X"6F",X"01",X"00",X"20",X"8D",X"E9",X"2C",X"04",X"A0",X"A9",X"4C",X"F7",
		X"2A",X"42",X"A9",X"94",X"D4",X"AA",X"44",X"52",X"D5",X"AA",X"AA",X"AA",X"EE",X"BE",X"DB",X"DA",
		X"6E",X"FF",X"DE",X"ED",X"2D",X"00",X"00",X"82",X"D0",X"BE",X"06",X"42",X"15",X"91",X"75",X"97",
		X"4A",X"A9",X"10",X"A9",X"56",X"55",X"15",X"80",X"ED",X"23",X"BF",X"56",X"BA",X"DB",X"D6",X"DB",
		X"FE",X"DF",X"DB",X"55",X"01",X"00",X"70",X"E8",X"D7",X"01",X"00",X"A5",X"F8",X"AF",X"41",X"0C",
		X"42",X"F5",X"AD",X"A9",X"0A",X"04",X"75",X"DD",X"D6",X"8A",X"54",X"BB",X"DD",X"5B",X"75",X"DF",
		X"FB",X"BF",X"DB",X"52",X"02",X"00",X"78",X"F8",X"4B",X"00",X"04",X"45",X"FD",X"95",X"A1",X"04",
		X"A4",X"3B",X"F5",X"AA",X"00",X"95",X"A8",X"FD",X"52",X"55",X"91",X"DE",X"DB",X"DE",X"DA",X"EE",
		X"FB",X"DF",X"B7",X"A6",X"34",X"00",X"80",X"81",X"3F",X"05",X"38",X"00",X"D5",X"47",X"4F",X"0B",
		X"30",X"A5",X"E8",X"97",X"A2",X"16",X"12",X"7C",X"D1",X"EA",X"43",X"AB",X"2E",X"FD",X"6E",X"ED",
		X"F7",X"DD",X"6F",X"57",X"55",X"01",X"00",X"10",X"F8",X"53",X"A1",X"02",X"88",X"5A",X"DC",X"B5",
		X"50",X"05",X"44",X"AD",X"EA",X"B6",X"A2",X"82",X"91",X"56",X"5F",X"5D",X"B5",X"F2",X"F5",X"DB",
		X"DF",X"F7",X"FE",X"B6",X"BD",X"12",X"00",X"00",X"A0",X"3E",X"5A",X"4A",X"80",X"48",X"4A",X"AF",
		X"5A",X"95",X"40",X"A2",X"A4",X"AD",X"6D",X"5D",X"A0",X"A2",X"A4",X"57",X"D7",X"36",X"ED",X"DD",
		X"FE",X"DD",X"FF",X"7B",X"77",X"BB",X"12",X"00",X"00",X"90",X"2E",X"AE",X"52",X"60",X"10",X"C5",
		X"55",X"AD",X"2A",X"52",X"48",X"54",X"A5",X"B5",X"AB",X"A8",X"22",X"51",X"AB",X"F5",X"B6",X"76",
		X"7B",X"EF",X"FB",X"FF",X"FE",X"6E",X"EB",X"25",X"80",X"00",X"00",X"07",X"5B",X"65",X"68",X"88",
		X"A2",X"49",X"2B",X"95",X"4A",X"28",X"A5",X"D2",X"AA",X"56",X"0B",X"35",X"2A",X"75",X"D1",X"BA",
		X"D5",X"6F",X"DF",X"6F",X"BF",X"BB",X"7B",X"6B",X"6B",X"05",X"08",X"00",X"62",X"A0",X"18",X"89",
		X"A3",X"54",X"2D",X"56",X"55",X"54",X"49",X"52",X"A5",X"54",X"55",X"55",X"B5",X"AA",X"AA",X"AA",
		X"4A",X"55",X"55",X"F5",X"DD",X"7D",X"DF",X"BD",X"BB",X"ED",X"DA",X"AE",X"0A",X"04",X"20",X"00",
		X"41",X"22",X"A5",X"AA",X"AA",X"5A",X"B5",X"A9",X"55",X"A5",X"94",X"24",X"8A",X"94",X"54",X"A9",
		X"AA",X"56",X"AB",X"AA",X"AA",X"7A",X"DD",X"EE",X"DD",X"FB",X"EE",X"77",X"77",X"5B",X"15",X"10",
		X"40",X"00",X"82",X"84",X"94",X"2A",X"55",X"AD",X"EA",X"6A",X"AB",X"2A",X"25",X"89",X"94",X"94",
		X"54",X"95",X"5A",X"D5",X"AA",X"EB",X"D6",X"EE",X"76",X"EF",X"DE",X"7B",X"BF",X"7B",X"5B",X"6B",
		X"01",X"0A",X"10",X"40",X"90",X"90",X"A2",X"4A",X"AB",X"5A",X"5D",X"AD",X"AA",X"54",X"51",X"A2",
		X"22",X"A5",X"4A",X"AA",X"AA",X"AA",X"5A",X"B7",X"75",X"B7",X"BD",X"BB",X"F7",X"DE",X"77",X"6F",
		X"6B",X"AB",X"80",X"00",X"01",X"04",X"09",X"49",X"2A",X"69",X"D5",X"AA",X"55",X"57",X"25",X"55",
		X"94",X"A4",X"28",X"A9",X"52",X"A9",X"4A",X"97",X"5E",X"5B",X"B7",X"BB",X"7D",X"7B",X"F7",X"BD",
		X"77",X"DB",X"D5",X"2A",X"20",X"40",X"00",X"42",X"22",X"92",X"4A",X"AA",X"6A",X"D5",X"AA",X"AB",
		X"94",X"2A",X"4A",X"2A",X"52",X"4A",X"55",X"52",X"55",X"AB",X"56",X"AF",X"DD",X"DE",X"BE",X"7B",
		X"F7",X"BD",X"BB",X"5B",X"6B",X"15",X"20",X"01",X"01",X"04",X"09",X"49",X"AA",X"54",X"D5",X"AA",
		X"D5",X"55",X"A5",X"4A",X"4A",X"52",X"54",X"52",X"A5",X"52",X"55",X"D5",X"BA",X"6E",X"BB",X"BB",
		X"77",X"EF",X"BD",X"F7",X"EE",X"6E",X"AB",X"55",X"40",X"80",X"00",X"42",X"44",X"94",X"54",X"AA",
		X"AA",X"55",X"AB",X"AB",X"AA",X"54",X"92",X"A4",X"A4",X"A4",X"4A",X"A9",X"4A",X"AB",X"6A",X"BD",
		X"DD",X"DD",X"7B",X"EF",X"DE",X"BB",X"77",X"B7",X"6D",X"55",X"01",X"02",X"04",X"20",X"44",X"24",
		X"A9",X"54",X"55",X"55",X"AD",X"DA",X"2A",X"A5",X"92",X"24",X"A5",X"94",X"2A",X"A9",X"54",X"55",
		X"DD",X"F5",X"EE",X"EE",X"BB",X"BB",X"77",X"6F",X"EF",X"76",X"6D",X"55",X"04",X"08",X"00",X"88",
		X"A0",X"48",X"A5",X"4A",X"55",X"AD",X"BA",X"B4",X"AA",X"52",X"49",X"4A",X"4A",X"52",X"A4",X"52",
		X"55",X"AB",X"5F",X"BF",X"BE",X"7D",X"BB",X"DB",X"B5",X"6B",X"AB",X"AD",X"5A",X"68",X"40",X"01",
		X"01",X"03",X"12",X"15",X"35",X"D9",X"AA",X"65",X"87",X"17",X"2D",X"1A",X"69",X"D0",X"A2",X"C5",
		X"CA",X"D5",X"CD",X"97",X"3E",X"7D",X"7C",X"F4",X"E2",X"E1",X"85",X"87",X"2E",X"AD",X"6E",X"A1",
		X"07",X"0E",X"0E",X"3C",X"70",X"B0",X"D0",X"85",X"8D",X"8E",X"4E",X"D5",X"4A",X"87",X"07",X"27",
		X"55",X"A9",X"D1",X"2A",X"1F",X"AF",X"BA",X"AE",X"8E",X"C7",X"96",X"36",X"9C",X"1C",X"A6",X"58",
		X"C5",X"D1",X"72",X"EA",X"EA",X"38",X"E3",X"8C",X"0B",X"0B",X"0E",X"0E",X"5C",X"58",X"E2",X"D0",
		X"E2",X"C4",X"35",X"76",X"F8",X"92",X"8F",X"E3",X"38",X"1C",X"F8",X"F0",X"C8",X"1C",X"75",X"F8",
		X"F0",X"E2",X"F1",X"F8",X"F0",X"98",X"0B",X"C7",X"C2",X"A3",X"E2",X"D0",X"B1",X"AA",X"AA",X"3A",
		X"3C",X"3C",X"3C",X"3C",X"0E",X"1F",X"3C",X"38",X"78",X"B8",X"78",X"3C",X"3C",X"3C",X"7C",X"78",
		X"8A",X"87",X"87",X"C3",X"85",X"0E",X"87",X"0F",X"0F",X"17",X"4F",X"95",X"B3",X"A6",X"86",X"2B",
		X"8E",X"0E",X"1E",X"0E",X"0F",X"9E",X"9A",X"72",X"6A",X"79",X"38",X"5E",X"78",X"D8",X"70",X"25",
		X"A7",X"3A",X"7C",X"F0",X"F0",X"E1",X"51",X"1E",X"1E",X"3C",X"1C",X"2B",X"0F",X"3E",X"0E",X"8F",
		X"C5",X"0B",X"1F",X"1E",X"3C",X"CA",X"91",X"17",X"8E",X"1E",X"F4",X"A8",X"E3",X"A1",X"87",X"2E",
		X"39",X"7A",X"F0",X"E0",X"C3",X"85",X"2F",X"3C",X"F4",X"58",X"1A",X"0F",X"3E",X"CC",X"29",X"65",
		X"07",X"1F",X"36",X"3C",X"D6",X"E1",X"98",X"0B",X"4F",X"36",X"0F",X"57",X"4E",X"9D",X"B2",X"0F",
		X"1E",X"8E",X"1E",X"53",X"E3",X"E4",X"E2",X"54",X"E3",X"B1",X"D0",X"C5",X"E4",X"51",X"55",X"A6",
		X"49",X"C3",X"E3",X"A8",X"94",X"A5",X"1A",X"B5",X"A8",X"0D",X"47",X"1B",X"1E",X"47",X"0F",X"8F",
		X"96",X"C6",X"5A",X"3A",X"2D",X"AD",X"5A",X"8E",X"8D",X"7C",X"28",X"8F",X"D4",X"25",X"69",X"43",
		X"3D",X"A8",X"4A",X"28",X"0B",X"B4",X"A0",X"56",X"51",X"2B",X"DA",X"49",X"AD",X"27",X"BD",X"6A",
		X"7D",X"6A",X"5F",X"F9",X"4D",X"F6",X"2A",X"BD",X"AA",X"DB",X"9B",X"F4",X"82",X"9A",X"24",X"55",
		X"95",X"BA",X"49",X"DD",X"2A",X"5F",X"75",X"57",X"6F",X"BD",X"DA",X"AD",X"7A",X"D5",X"AA",X"55",
		X"D8",X"48",X"4A",X"02",X"15",X"24",X"22",X"91",X"04",X"20",X"02",X"40",X"20",X"20",X"82",X"44",
		X"24",X"29",X"55",X"55",X"B5",X"D6",X"B6",X"B5",X"6D",X"DB",X"B6",X"ED",X"EE",X"EE",X"FB",X"BE",
		X"EF",X"F7",X"DE",X"BB",X"BB",X"BB",X"DB",X"EE",X"B6",X"6D",X"AB",X"2A",X"91",X"88",X"24",X"94",
		X"92",X"AA",X"54",X"B5",X"AA",X"AB",X"AA",X"4A",X"89",X"88",X"10",X"22",X"49",X"52",X"55",X"AD",
		X"F6",X"B6",X"AD",X"6D",X"B5",X"AA",X"2A",X"55",X"01",X"10",X"00",X"80",X"20",X"90",X"24",X"55",
		X"AA",X"AA",X"55",X"DB",X"6A",X"AD",X"AA",X"52",X"29",X"22",X"4A",X"52",X"D5",X"77",X"7F",X"7F",
		X"EF",X"6F",X"6F",X"77",X"BB",X"6D",X"17",X"29",X"20",X"00",X"24",X"50",X"A9",X"2A",X"B5",X"D5",
		X"AD",X"6E",X"B5",X"D5",X"AA",X"AA",X"A4",X"24",X"45",X"54",X"52",X"D5",X"BE",X"7F",X"7F",X"DF",
		X"DF",X"BD",X"BB",X"77",X"77",X"13",X"25",X"00",X"00",X"11",X"28",X"A9",X"92",X"5A",X"D5",X"D2",
		X"AB",X"B6",X"AA",X"8A",X"4A",X"92",X"48",X"21",X"49",X"2A",X"D5",X"DE",X"EF",X"FD",X"FD",X"BE",
		X"EF",X"DE",X"DD",X"5B",X"85",X"08",X"00",X"80",X"04",X"4A",X"54",X"49",X"AD",X"5A",X"D5",X"AD",
		X"55",X"B5",X"28",X"49",X"49",X"92",X"48",X"89",X"4A",X"AD",X"ED",X"DF",X"DF",X"EF",X"F7",X"7B",
		X"EF",X"DE",X"DD",X"8A",X"88",X"00",X"00",X"12",X"28",X"51",X"95",X"AA",X"DA",X"AA",X"6B",X"5B",
		X"55",X"A5",X"24",X"92",X"24",X"14",X"89",X"B4",X"B2",X"BF",X"7D",X"7F",X"FB",X"DF",X"EF",X"DB",
		X"DF",X"BD",X"05",X"1C",X"00",X"00",X"49",X"82",X"16",X"D8",X"50",X"AB",X"AD",X"5E",X"BC",X"50",
		X"45",X"25",X"95",X"54",X"A5",X"4A",X"55",X"F5",X"BA",X"DB",X"BB",X"EF",X"FE",X"FE",X"FE",X"FA",
		X"EB",X"AF",X"06",X"07",X"08",X"C0",X"80",X"05",X"85",X"0A",X"3D",X"F8",X"E1",X"8B",X"8E",X"54",
		X"54",X"54",X"A1",X"83",X"0E",X"6D",X"B4",X"E9",X"EA",X"D6",X"5D",X"6F",X"7D",X"FB",X"ED",X"FB",
		X"F6",X"5E",X"17",X"1C",X"10",X"C0",X"80",X"03",X"16",X"2C",X"5C",X"F4",X"F0",X"85",X"17",X"1D",
		X"AA",X"A8",X"A4",X"52",X"93",X"3C",X"F8",X"E1",X"43",X"1F",X"5F",X"EE",X"DA",X"76",X"FD",X"D5",
		X"AF",X"AF",X"D5",X"C1",X"01",X"01",X"1C",X"30",X"B0",X"50",X"C3",X"4A",X"4B",X"97",X"BC",X"E8",
		X"50",X"45",X"4A",X"4A",X"55",X"5A",X"F4",X"E8",X"45",X"4F",X"37",X"DD",X"DA",X"6D",X"EF",X"F6",
		X"FB",X"B7",X"77",X"D7",X"82",X"03",X"02",X"18",X"30",X"D0",X"82",X"A3",X"AA",X"54",X"4B",X"5B",
		X"3A",X"52",X"A1",X"44",X"2A",X"A5",X"AA",X"56",X"7A",X"F8",X"E0",X"C3",X"87",X"2F",X"AF",X"76",
		X"BB",X"BB",X"BF",X"BE",X"F5",X"52",X"38",X"10",X"C0",X"80",X"02",X"17",X"5A",X"54",X"4B",X"AD",
		X"74",X"D1",X"49",X"15",X"2A",X"A9",X"A4",X"AA",X"5A",X"AD",X"AD",X"B6",X"6C",X"71",X"D5",X"D5",
		X"EB",X"EE",X"DE",X"FB",X"BE",X"7B",X"7B",X"D5",X"E0",X"00",X"00",X"03",X"12",X"1C",X"AA",X"51",
		X"2D",X"D5",X"68",X"A5",X"A3",X"2A",X"2A",X"51",X"49",X"95",X"6A",X"B5",X"3A",X"7C",X"F8",X"E0",
		X"C3",X"8B",X"5E",X"5D",X"BB",X"BB",X"BB",X"BD",X"ED",X"D6",X"AA",X"70",X"10",X"80",X"01",X"11",
		X"0E",X"75",X"58",X"8B",X"35",X"5C",X"D2",X"A1",X"26",X"96",X"A8",X"A4",X"2A",X"AB",X"5A",X"1D",
		X"1F",X"5E",X"78",X"E8",X"62",X"57",X"57",X"77",X"BB",X"BB",X"B7",X"B7",X"5E",X"B5",X"82",X"83",
		X"01",X"0C",X"48",X"70",X"A8",X"A3",X"3A",X"5C",X"D1",X"45",X"8B",X"5A",X"68",X"51",X"95",X"AA",
		X"B4",X"EA",X"3A",X"BC",X"78",X"E1",X"45",X"17",X"37",X"DD",X"BA",X"DB",X"DB",X"BD",X"6E",X"6D",
		X"D5",X"02",X"1E",X"0C",X"60",X"20",X"82",X"C3",X"1A",X"EB",X"B0",X"15",X"17",X"3A",X"D4",X"A2",
		X"4A",X"56",X"AA",X"D2",X"AA",X"2E",X"8F",X"AB",X"5A",X"5C",X"74",X"A9",X"6B",X"B7",X"7B",X"F7",
		X"ED",X"6D",X"B7",X"56",X"4D",X"05",X"07",X"02",X"38",X"50",X"C0",X"51",X"47",X"75",X"68",X"43",
		X"8B",X"1C",X"69",X"A1",X"25",X"2B",X"B5",X"D4",X"AA",X"9B",X"7C",X"78",X"F0",X"C1",X"0B",X"2F",
		X"BD",X"DA",X"B6",X"B7",X"BD",X"F6",X"6A",X"CB",X"4A",X"05",X"0E",X"0A",X"70",X"60",X"C1",X"45",
		X"1D",X"B3",X"52",X"0B",X"17",X"3A",X"D4",X"A4",X"4A",X"55",X"6A",X"A5",X"55",X"B7",X"F0",X"E0",
		X"C1",X"07",X"0F",X"1F",X"DE",X"74",X"6B",X"B7",X"BD",X"7A",X"D5",X"A5",X"95",X"0A",X"1C",X"28",
		X"E0",X"C0",X"82",X"4B",X"B5",X"54",X"53",X"95",X"54",X"D1",X"48",X"93",X"2A",X"55",X"55",X"55",
		X"BB",X"EA",X"F2",X"52",X"87",X"2E",X"BA",X"E8",X"EA",X"B6",X"BB",X"7D",X"7B",X"D7",X"AB",X"5B",
		X"6A",X"A1",X"02",X"0D",X"04",X"70",X"60",X"85",X"53",X"56",X"AA",X"A9",X"4A",X"96",X"58",X"51",
		X"A5",X"2A",X"55",X"D5",X"AA",X"AB",X"6E",X"F8",X"F0",X"C0",X"87",X"07",X"1F",X"BD",X"BA",X"B5",
		X"DB",X"76",X"ED",X"D5",X"A6",X"16",X"1A",X"A2",X"81",X"01",X"2E",X"58",X"E8",X"A4",X"96",X"AA",
		X"54",X"45",X"15",X"2D",X"B2",X"A4",X"4A",X"2D",X"B5",X"AA",X"53",X"55",X"55",X"95",X"AA",X"AA",
		X"5A",X"BD",X"BD",X"BB",X"F7",X"DE",X"DE",X"6E",X"5B",X"AB",X"2A",X"94",X"10",X"02",X"43",X"18",
		X"54",X"D1",X"52",X"4D",X"55",X"AA",X"92",X"4A",X"AA",X"54",X"A9",X"4A",X"55",X"B5",X"EA",X"55",
		X"97",X"96",X"B4",X"54",X"55",X"55",X"7B",X"7D",X"7B",X"BB",X"77",X"B7",X"DB",X"B6",X"D5",X"AA",
		X"22",X"09",X"09",X"02",X"09",X"2A",X"A4",X"52",X"A5",X"AA",X"54",X"A9",X"92",X"4A",X"AA",X"54",
		X"A9",X"4A",X"55",X"D5",X"6A",X"5D",X"2D",X"55",X"55",X"55",X"55",X"BD",X"DB",X"BD",X"BB",X"77",
		X"B7",X"BB",X"6E",X"6B",X"AD",X"4A",X"A1",X"88",X"08",X"41",X"84",X"28",X"52",X"51",X"A5",X"AA",
		X"54",X"A9",X"52",X"2A",X"55",X"AA",X"54",X"55",X"55",X"AD",X"55",X"57",X"57",X"AD",X"54",X"D5",
		X"A5",X"EB",X"B6",X"BB",X"BB",X"BB",X"BB",X"DD",X"B6",X"6D",X"AD",X"AA",X"82",X"82",X"82",X"24",
		X"28",X"A4",X"48",X"49",X"95",X"AA",X"52",X"2A",X"55",X"52",X"49",X"29",X"95",X"AA",X"54",X"55",
		X"B5",X"EA",X"A5",X"AA",X"2A",X"55",X"B5",X"EA",X"EB",X"6E",X"6F",X"77",X"B7",X"BB",X"DD",X"B6",
		X"AD",X"56",X"55",X"A0",X"88",X"82",X"12",X"92",X"28",X"91",X"4A",X"AA",X"54",X"A5",X"4A",X"95",
		X"54",X"52",X"25",X"55",X"AA",X"AA",X"AA",X"D5",X"AA",X"4A",X"8B",X"96",X"BA",X"6A",X"D5",X"D7",
		X"DB",X"DE",X"EE",X"B6",X"BB",X"ED",X"D6",X"D6",X"AA",X"24",X"28",X"22",X"41",X"22",X"8A",X"24",
		X"29",X"29",X"55",X"AA",X"54",X"29",X"95",X"52",X"52",X"A5",X"AA",X"AA",X"6A",X"AD",X"3A",X"55",
		X"A5",X"95",X"56",X"AD",X"EA",X"DB",X"DB",X"DD",X"6E",X"BB",X"DB",X"5D",X"AF",X"6D",X"B5",X"8A",
		X"82",X"22",X"14",X"92",X"90",X"44",X"92",X"A4",X"94",X"AA",X"54",X"AA",X"94",X"4A",X"A5",X"54",
		X"AA",X"AA",X"AA",X"AD",X"7A",X"A9",X"AA",X"AA",X"AA",X"7A",X"DD",X"DA",X"ED",X"6D",X"77",X"BB",
		X"DB",X"DD",X"76",X"6D",X"6B",X"2B",X"55",X"50",X"88",X"08",X"11",X"12",X"91",X"24",X"25",X"55",
		X"AA",X"94",X"4A",X"29",X"A5",X"A4",X"4A",X"55",X"55",X"55",X"5D",X"6C",X"F1",X"A2",X"57",X"5B",
		X"5D",X"BD",X"B5",X"DB",X"6E",X"BB",X"BB",X"DD",X"6E",X"BB",X"B5",X"AA",X"22",X"21",X"09",X"22",
		X"42",X"84",X"12",X"95",X"54",X"A9",X"4A",X"A5",X"94",X"52",X"4A",X"2A",X"55",X"A9",X"AA",X"AA",
		X"96",X"0E",X"5F",X"78",X"F1",X"E2",X"55",X"57",X"5D",X"ED",X"DA",X"6E",X"77",X"DB",X"6D",X"5B",
		X"5B",X"55",X"89",X"24",X"A2",X"40",X"42",X"0A",X"2A",X"4A",X"A9",X"52",X"95",X"AA",X"94",X"2A",
		X"55",X"52",X"A5",X"AA",X"AA",X"AA",X"D5",X"6E",X"8B",X"0F",X"1F",X"7C",X"F8",X"F0",X"A5",X"97",
		X"AE",X"B5",X"6D",X"BB",X"BA",X"DA",X"6A",X"4B",X"0B",X"25",X"92",X"44",X"0A",X"29",X"A2",X"48",
		X"92",X"94",X"52",X"A9",X"52",X"A9",X"52",X"A5",X"4A",X"55",X"55",X"B5",X"6A",X"D5",X"AD",X"55",
		X"5B",X"AA",X"EA",X"AB",X"DB",X"B6",X"ED",X"ED",X"6D",X"77",X"7B",X"BB",X"6D",X"6B",X"AB",X"AA",
		X"22",X"44",X"82",X"12",X"2A",X"54",X"A2",X"44",X"89",X"8A",X"54",X"A9",X"94",X"52",X"4A",X"29",
		X"55",X"55",X"55",X"AB",X"55",X"55",X"55",X"D5",X"5B",X"5D",X"74",X"E9",X"EA",X"55",X"57",X"B7",
		X"B6",X"76",X"ED",X"DA",X"D5",X"AD",X"AD",X"AE",X"B6",X"6A",X"55",X"22",X"89",X"48",X"48",X"22",
		X"45",X"2A",X"54",X"51",X"49",X"2A",X"29",X"A9",X"24",X"A5",X"2A",X"AA",X"AA",X"6A",X"B5",X"D7",
		X"B6",X"6D",X"DD",X"DA",X"B6",X"5B",X"DB",X"5A",X"AB",X"AA",X"A2",X"52",X"85",X"0A",X"55",X"54",
		X"A5",X"42",X"0B",X"55",X"54",X"A9",X"A2",X"4A",X"A5",X"AA",X"AA",X"BA",X"AA",X"6B",X"5B",X"6D",
		X"5B",X"6B",X"AB",X"5B",X"BB",X"B6",X"AD",X"AE",X"B6",X"6A",X"A9",X"24",X"49",X"91",X"90",X"22",
		X"49",X"92",X"12",X"95",X"94",X"92",X"92",X"44",X"15",X"5A",X"AA",X"AA",X"AA",X"D6",X"56",X"DF",
		X"7A",X"B5",X"AD",X"AD",X"B6",X"B5",X"6A",X"AB",X"37",X"F9",X"F8",X"82",X"83",X"2A",X"AA",X"A8",
		X"A2",X"A2",X"2A",X"55",X"69",X"55",X"55",X"55",X"A5",X"2A",X"55",X"AA",X"AA",X"D6",X"7A",X"DB",
		X"5E",X"7B",X"B5",X"AD",X"6E",X"B5",X"AD",X"B6",X"5A",X"B5",X"5A",X"4A",X"49",X"0A",X"91",X"08",
		X"09",X"52",X"48",X"49",X"92",X"8A",X"AA",X"54",X"55",X"55",X"55",X"AB",X"AA",X"55",X"55",X"55",
		X"5F",X"ED",X"6A",X"D5",X"AB",X"AE",X"BA",X"EA",X"AA",X"55",X"2D",X"95",X"AA",X"54",X"55",X"A9",
		X"4A",X"2A",X"B4",X"50",X"A1",X"8A",X"2A",X"2A",X"AA",X"A2",X"AA",X"2A",X"55",X"55",X"B5",X"6A",
		X"55",X"BD",X"6A",X"D7",X"B6",X"55",X"57",X"B5",X"B5",X"B5",X"9A",X"AA",X"52",X"2B",X"55",X"51",
		X"AD",X"A8",X"8E",X"AA",X"42",X"2B",X"AA",X"A2",X"94",X"50",X"89",X"92",X"A8",X"A4",X"54",X"A5",
		X"55",X"DB",X"DB",X"6E",X"ED",X"56",X"57",X"DB",X"B6",X"BA",X"DA",X"D6",X"6E",X"B5",X"D5",X"AA",
		X"AB",X"52",X"A8",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"2A",X"00",X"00",X"00",X"F8",X"5F",
		X"EF",X"B7",X"6E",X"5D",X"6B",X"55",X"00",X"50",X"AB",X"8A",X"D4",X"BD",X"9B",X"AA",X"6D",X"21",
		X"ED",X"FF",X"DD",X"FD",X"DF",X"F7",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"00",X"D0",X"76",
		X"89",X"AD",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"81",X"20",X"44",X"44",X"C5",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"0F",X"C4",X"FF",X"DF",X"37",X"04",
		X"25",X"48",X"FD",X"5F",X"00",X"00",X"90",X"D2",X"56",X"03",X"08",X"ED",X"DB",X"A5",X"AB",X"5F",
		X"00",X"00",X"F8",X"FF",X"07",X"00",X"00",X"00",X"F8",X"FF",X"01",X"00",X"00",X"A0",X"FF",X"1F",
		X"00",X"80",X"FE",X"FD",X"7F",X"03",X"00",X"FA",X"FF",X"2F",X"A5",X"54",X"FF",X"FF",X"7F",X"A9",
		X"FF",X"FF",X"FF",X"0F",X"00",X"C0",X"FF",X"7F",X"04",X"00",X"00",X"FD",X"FF",X"07",X"00",X"B6",
		X"BD",X"FF",X"3F",X"00",X"F0",X"FF",X"FF",X"BF",X"09",X"40",X"FF",X"FF",X"4D",X"20",X"A9",X"FF",
		X"FF",X"15",X"44",X"FD",X"FF",X"FF",X"37",X"00",X"00",X"FC",X"FF",X"63",X"10",X"00",X"D0",X"FF",
		X"1F",X"00",X"A9",X"A8",X"FF",X"FF",X"02",X"40",X"FB",X"BD",X"FF",X"95",X"00",X"D5",X"FE",X"7F",
		X"95",X"40",X"F4",X"FF",X"DF",X"2A",X"55",X"FB",X"FF",X"FB",X"6F",X"01",X"00",X"00",X"FE",X"5B",
		X"09",X"00",X"00",X"D0",X"BF",X"AB",X"02",X"00",X"F0",X"FE",X"D6",X"55",X"09",X"A0",X"FE",X"FF",
		X"5D",X"2B",X"44",X"F5",X"FF",X"6E",X"B5",X"DD",X"FB",X"DF",X"6F",X"77",X"FF",X"FF",X"FF",X"5F",
		X"00",X"00",X"20",X"FD",X"FE",X"04",X"00",X"00",X"90",X"EE",X"BE",X"12",X"00",X"10",X"25",X"5B",
		X"B7",X"55",X"48",X"48",X"C9",X"AA",X"6E",X"57",X"12",X"94",X"A4",X"EA",X"FF",X"BF",X"AD",X"AD",
		X"D6",X"FE",X"FF",X"FF",X"23",X"00",X"00",X"00",X"DA",X"77",X"AD",X"2A",X"00",X"90",X"54",X"B7",
		X"7F",X"37",X"25",X"51",X"69",X"6D",X"DB",X"6E",X"55",X"DB",X"B5",X"2A",X"25",X"55",X"7B",X"FF",
		X"BB",X"B5",X"76",X"BB",X"BB",X"5B",X"2B",X"D5",X"FD",X"4D",X"00",X"00",X"00",X"00",X"48",X"A9",
		X"AA",X"84",X"20",X"91",X"28",X"55",X"55",X"AA",X"AA",X"A5",X"44",X"49",X"95",X"5A",X"BB",X"B5",
		X"AA",X"AA",X"B2",X"99",X"66",X"CE",X"DC",X"DD",X"D9",X"DE",X"CE",X"14",X"69",X"62",X"DF",X"0A",
		X"02",X"00",X"00",X"24",X"11",X"24",X"51",X"C6",X"AA",X"D6",X"98",X"A9",X"DE",X"7A",X"77",X"CE",
		X"8C",X"39",X"7B",X"33",X"67",X"CE",X"6C",X"77",X"67",X"D7",X"CC",X"EC",X"9C",X"BD",X"6D",X"4C",
		X"96",X"6C",X"67",X"CE",X"10",X"88",X"11",X"33",X"26",X"22",X"00",X"40",X"12",X"22",X"26",X"62",
		X"C6",X"A4",X"64",X"CE",X"CC",X"9D",X"1D",X"1B",X"39",X"33",X"B7",X"56",X"29",X"D9",X"9D",X"DD",
		X"CD",X"6D",X"D5",X"5C",X"33",X"73",X"CE",X"6E",X"96",X"98",X"C4",X"9C",X"99",X"35",X"22",X"22",
		X"64",X"26",X"04",X"21",X"26",X"62",X"8A",X"19",X"99",X"31",X"53",X"76",X"EE",X"CC",X"DC",X"99",
		X"39",X"73",X"76",X"B7",X"97",X"71",X"56",X"99",X"BD",X"1A",X"63",X"32",X"49",X"4A",X"84",X"88",
		X"09",X"11",X"89",X"92",X"8C",X"18",X"73",X"66",X"6C",X"6D",X"A6",X"9D",X"CD",X"98",X"63",X"CE",
		X"DC",X"9C",X"55",X"31",X"76",X"E6",X"66",X"92",X"19",X"93",X"C4",X"24",X"A9",X"64",X"66",X"2C",
		X"21",X"C5",X"D0",X"CC",X"99",X"19",X"73",X"CC",X"98",X"99",X"35",X"66",X"CE",X"98",X"67",X"8C",
		X"99",X"94",X"59",X"73",X"CE",X"60",X"CA",X"9C",X"31",X"CE",X"18",X"CB",X"39",X"63",X"66",X"CC",
		X"33",X"E7",X"8C",X"74",X"C6",X"38",X"D7",X"26",X"B3",X"9D",X"33",X"8F",X"33",X"6B",X"35",X"C9",
		X"31",X"67",X"8C",X"99",X"09",X"B3",X"8C",X"8D",X"CC",X"68",X"AC",X"39",X"66",X"CC",X"31",X"E7",
		X"19",X"D7",X"98",X"EB",X"9C",X"66",X"9C",X"B9",X"E6",X"D6",X"CA",X"19",X"93",X"19",X"23",X"84",
		X"88",X"08",X"53",X"94",X"2A",X"A6",X"D6",X"D8",X"9A",X"DA",X"33",X"EF",X"AC",X"DB",X"39",X"D7",
		X"5D",X"E7",X"9E",X"73",X"CF",X"39",X"AF",X"11",X"84",X"00",X"A0",X"10",X"D5",X"4A",X"55",X"25",
		X"55",X"4A",X"55",X"AD",X"BA",X"56",X"15",X"A3",X"94",X"54",X"5D",X"FD",X"7A",X"F7",X"F6",X"B6",
		X"EB",X"DD",X"77",X"DF",X"5D",X"B7",X"0A",X"01",X"00",X"00",X"45",X"4A",X"B5",X"54",X"A5",X"A4",
		X"92",X"AA",X"B5",X"6E",X"AD",X"AA",X"22",X"A5",X"52",X"BD",X"7D",X"B7",X"AD",X"B5",X"75",X"F7",
		X"DE",X"F7",X"DD",X"7D",X"7F",X"6F",X"15",X"00",X"00",X"00",X"A0",X"AA",X"95",X"56",X"44",X"14",
		X"94",X"6A",X"AD",X"57",X"AB",X"2A",X"AA",X"54",X"A3",X"DB",X"B6",X"6F",X"DD",X"5A",X"6D",X"DB",
		X"FB",X"FE",X"BD",X"FB",X"EE",X"7B",X"DF",X"64",X"01",X"00",X"00",X"00",X"5A",X"B5",X"D2",X"04",
		X"48",X"82",X"5A",X"B5",X"77",X"55",X"2B",X"92",X"2A",X"55",X"D9",X"ED",X"F6",X"B6",X"AD",X"AE",
		X"BA",X"DB",X"FB",X"EF",X"DF",X"F7",X"BD",X"5B",X"54",X"00",X"00",X"00",X"20",X"6C",X"AA",X"4A",
		X"81",X"44",X"48",X"5A",X"75",X"D7",X"D6",X"4A",X"29",X"A9",X"AA",X"FC",X"BA",X"FB",X"D6",X"AE",
		X"EA",X"6A",X"F7",X"F7",X"FD",X"FB",X"BD",X"EF",X"DE",X"92",X"01",X"00",X"00",X"00",X"42",X"97",
		X"AA",X"22",X"88",X"02",X"95",X"B4",X"B5",X"B5",X"56",X"54",X"52",X"AA",X"74",X"DB",X"FB",X"AE",
		X"5B",X"A5",X"55",X"FB",X"FB",X"FF",X"DE",X"DF",X"EE",X"BB",X"AD",X"64",X"00",X"00",X"00",X"00",
		X"D1",X"25",X"B5",X"40",X"22",X"48",X"AA",X"EA",X"56",X"5B",X"55",X"52",X"45",X"BA",X"EA",X"B7",
		X"BB",X"B7",X"AA",X"95",X"76",X"F7",X"EF",X"BF",X"BF",X"DD",X"6F",X"7B",X"43",X"05",X"00",X"00",
		X"00",X"A0",X"5A",X"D2",X"0A",X"24",X"88",X"A4",X"AA",X"B6",X"DA",X"96",X"4A",X"25",X"D2",X"A5",
		X"FE",X"F6",X"BB",X"AD",X"B6",X"EA",X"5E",X"FF",X"DF",X"7F",X"F7",X"BD",X"BB",X"95",X"0A",X"00",
		X"00",X"00",X"80",X"AA",X"4A",X"2E",X"20",X"09",X"94",X"94",X"B6",X"55",X"B7",X"A8",X"2A",X"D2",
		X"4A",X"FD",X"B5",X"BF",X"75",X"B5",X"AA",X"BB",X"FD",X"DF",X"7F",X"F7",X"DE",X"6E",X"AB",X"92",
		X"00",X"00",X"00",X"00",X"48",X"A5",X"6A",X"81",X"0A",X"50",X"45",X"DA",X"AA",X"B6",X"55",X"AD",
		X"A0",X"27",X"DA",X"AB",X"BF",X"EB",X"AD",X"55",X"5B",X"DB",X"DF",X"FF",X"F5",X"5E",X"DB",X"D5",
		X"2A",X"05",X"00",X"00",X"00",X"80",X"88",X"AC",X"4A",X"AA",X"82",X"2A",X"A1",X"95",X"6C",X"A5",
		X"6E",X"55",X"B5",X"95",X"7E",X"F5",X"AF",X"DE",X"D6",X"56",X"DB",X"DA",X"ED",X"BE",X"DD",X"56",
		X"5B",X"55",X"55",X"14",X"00",X"00",X"00",X"00",X"0A",X"A4",X"12",X"6A",X"51",X"B5",X"D4",X"AA",
		X"DA",X"AA",X"5A",X"95",X"AA",X"AA",X"AA",X"B4",X"AB",X"DD",X"DA",X"B5",X"6A",X"AD",X"6E",X"DB",
		X"DD",X"76",X"AB",X"D5",X"4A",X"25",X"49",X"22",X"04",X"04",X"00",X"20",X"08",X"42",X"24",X"52",
		X"A9",X"AA",X"D5",X"6E",X"DB",X"AD",X"56",X"AB",X"2A",X"AA",X"AA",X"AA",X"AE",X"DD",X"BA",X"6D",
		X"77",X"77",X"B7",X"DB",X"5A",X"AD",X"2A",X"4A",X"92",X"14",X"91",X"20",X"02",X"10",X"00",X"02",
		X"42",X"48",X"22",X"95",X"AA",X"6A",X"AD",X"5B",X"5B",X"5B",X"6B",X"B5",X"AA",X"5A",X"55",X"5B",
		X"ED",X"6E",X"EF",X"BD",X"BB",X"DB",X"6E",X"D5",X"AA",X"AA",X"AA",X"94",X"2A",X"25",X"21",X"02",
		X"02",X"08",X"40",X"10",X"22",X"92",X"52",X"AA",X"AA",X"5A",X"EB",X"DA",X"D6",X"56",X"AB",X"AA",
		X"52",X"AA",X"6A",X"BD",X"BB",X"F7",X"EE",X"76",X"BB",X"AD",X"B5",X"5A",X"55",X"AD",X"2A",X"49",
		X"49",X"44",X"08",X"02",X"10",X"40",X"10",X"12",X"29",X"A5",X"AA",X"AA",X"B6",X"6B",X"DB",X"AE",
		X"AD",X"AA",X"AA",X"14",X"E0",X"47",X"FF",X"F5",X"AD",X"57",X"5D",X"AB",X"B6",X"5A",X"55",X"AB",
		X"A5",X"A2",X"92",X"22",X"84",X"00",X"01",X"02",X"22",X"44",X"92",X"4A",X"55",X"D5",X"5A",X"DB",
		X"6A",X"AB",X"AA",X"55",X"55",X"DD",X"DA",X"DD",X"FB",X"EE",X"DD",X"6D",X"DB",X"6A",X"D5",X"AA",
		X"5A",X"55",X"2A",X"25",X"49",X"04",X"21",X"08",X"10",X"10",X"22",X"49",X"4A",X"55",X"55",X"EB",
		X"6D",X"B7",X"6D",X"6B",X"AB",X"B5",X"D6",X"B6",X"ED",X"76",X"B7",X"ED",X"D6",X"B6",X"5A",X"55",
		X"15",X"AA",X"94",X"52",X"4A",X"A4",X"88",X"88",X"48",X"44",X"24",X"12",X"29",X"49",X"A9",X"4A",
		X"55",X"AD",X"56",X"F5",X"5A",X"6B",X"AB",X"6D",X"6B",X"DB",X"D6",X"B6",X"D6",X"B6",X"56",X"2B",
		X"4A",X"92",X"48",X"29",X"4A",X"49",X"A4",X"24",X"4A",X"24",X"09",X"25",X"92",X"A4",X"24",X"A9",
		X"52",X"95",X"AA",X"6A",X"AB",X"D5",X"AA",X"AA",X"EA",X"B5",X"DB",X"B6",X"DB",X"DA",X"AE",X"AA",
		X"AB",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"A8",X"2A",X"29",X"A5",X"28",X"55",
		X"55",X"55",X"AB",X"5A",X"55",X"55",X"AB",X"AA",X"AA",X"4A",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"92",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"4A",X"55",X"55",X"55",X"55",X"AB",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"56",X"55",X"55",X"55",X"95",X"AA",X"AA",X"B5",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"A5",
		X"AA",X"AA",X"AA",X"52",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"6D",X"55",X"55",X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"B5",X"5A",X"55",X"55",
		X"55",X"55",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"24",X"51",X"94",X"14",X"95",X"4A",X"55",X"55",
		X"55",X"55",X"B5",X"AA",X"AA",X"D5",X"AA",X"2A",X"00",X"00",X"E0",X"81",X"FF",X"FF",X"FF",X"F5",
		X"2F",X"E0",X"03",X"7E",X"D8",X"6F",X"D1",X"07",X"5E",X"90",X"16",X"F0",X"C1",X"5B",X"AA",X"8B",
		X"FA",X"F4",X"DF",X"FF",X"FD",X"07",X"00",X"00",X"00",X"FE",X"E1",X"0F",X"1C",X"00",X"08",X"FF",
		X"F9",X"AF",X"0F",X"20",X"05",X"FF",X"FE",X"FF",X"2D",X"78",X"C0",X"E7",X"FF",X"DD",X"97",X"5E",
		X"BE",X"7F",X"FF",X"FF",X"0F",X"02",X"00",X"80",X"FA",X"FA",X"22",X"00",X"00",X"20",X"DB",X"DF",
		X"9B",X"14",X"80",X"48",X"FD",X"FD",X"DF",X"5A",X"22",X"C4",X"BA",X"FF",X"BD",X"AB",X"55",X"B7",
		X"FF",X"FF",X"FF",X"7F",X"22",X"00",X"00",X"E5",X"EB",X"D3",X"02",X"00",X"00",X"A9",X"B7",X"5D",
		X"11",X"00",X"80",X"64",X"BD",X"D7",X"95",X"08",X"10",X"C9",X"F2",X"D5",X"C3",X"82",X"A2",X"AA",
		X"EF",X"BF",X"DF",X"FF",X"FB",X"82",X"00",X"00",X"D0",X"B4",X"D7",X"56",X"80",X"00",X"44",X"ED",
		X"FE",X"DD",X"4A",X"88",X"90",X"EA",X"FE",X"F7",X"B6",X"A4",X"A4",X"D6",X"F2",X"C3",X"87",X"0E",
		X"EB",X"DA",X"DF",X"BF",X"7F",X"FF",X"B6",X"14",X"20",X"00",X"20",X"AA",X"6A",X"A9",X"08",X"10",
		X"44",X"B2",X"DA",X"75",X"55",X"44",X"08",X"51",X"75",X"DF",X"EF",X"B6",X"52",X"89",X"14",X"0F",
		X"3E",X"FC",X"BC",X"D5",X"9E",X"7E",X"FF",X"FF",X"BF",X"0F",X"15",X"00",X"00",X"A4",X"AA",X"AE",
		X"34",X"82",X"80",X"44",X"AA",X"B6",X"5A",X"95",X"24",X"4A",X"AA",X"D5",X"B7",X"DD",X"6A",X"55",
		X"2B",X"51",X"24",X"71",X"E9",X"BB",X"7B",X"7B",X"DB",X"EE",X"7E",X"FF",X"FF",X"5A",X"08",X"00",
		X"00",X"20",X"A9",X"D2",X"52",X"91",X"20",X"42",X"94",X"AC",X"B5",X"B6",X"AA",X"24",X"25",X"D5",
		X"7A",X"B7",X"B7",X"6D",X"69",X"41",X"85",X"4B",X"BF",X"BF",X"FD",X"7A",X"EB",X"EB",X"6F",X"7F",
		X"5F",X"8D",X"04",X"00",X"00",X"22",X"28",X"49",X"A9",X"92",X"92",X"24",X"24",X"49",X"A9",X"5A",
		X"BB",X"B6",X"AA",X"4A",X"AA",X"DB",X"DD",X"D6",X"A3",X"8B",X"4B",X"AF",X"BF",X"7F",X"BF",X"6F",
		X"EF",X"F6",X"7D",X"ED",X"A4",X"02",X"02",X"00",X"08",X"24",X"54",X"52",X"A5",X"92",X"8A",X"94",
		X"94",X"54",X"A9",X"6A",X"B5",X"56",X"55",X"45",X"95",X"4A",X"AB",X"AE",X"7B",X"FD",X"F6",X"F7",
		X"FD",X"F7",X"BE",X"6F",X"B7",X"AA",X"40",X"00",X"00",X"02",X"04",X"25",X"55",X"AA",X"AA",X"A4",
		X"A2",X"24",X"95",X"AA",X"AA",X"55",X"4B",X"4B",X"D7",X"D5",X"DB",X"EE",X"6E",X"BB",X"FB",X"DE",
		X"EF",X"EF",X"77",X"B7",X"55",X"8B",X"02",X"01",X"00",X"00",X"10",X"22",X"49",X"A5",X"AA",X"55",
		X"55",X"4A",X"49",X"4A",X"4A",X"55",X"AD",X"AE",X"D7",X"D5",X"D7",X"EB",X"BB",X"EF",X"EE",X"B6",
		X"6D",X"D7",X"6D",X"AF",X"96",X"0A",X"04",X"00",X"00",X"40",X"50",X"92",X"AA",X"56",X"55",X"55",
		X"A5",X"52",X"52",X"52",X"A9",X"52",X"D5",X"6B",X"DF",X"FB",X"BE",X"77",X"77",X"BB",X"6E",X"DD",
		X"B6",X"56",X"25",X"02",X"01",X"00",X"00",X"09",X"49",X"AA",X"AA",X"AA",X"AA",X"AA",X"52",X"49",
		X"22",X"49",X"4A",X"AA",X"BD",X"EF",X"FB",X"7D",X"F7",X"DE",X"6E",X"DB",X"56",X"AD",X"14",X"89",
		X"40",X"20",X"40",X"08",X"89",X"54",X"4A",X"55",X"55",X"55",X"55",X"55",X"55",X"52",X"4A",X"4A",
		X"55",X"B5",X"F7",X"EE",X"BB",X"BB",X"DB",X"B6",X"D6",X"AA",X"56",X"D5",X"AA",X"92",X"44",X"22",
		X"84",X"88",X"44",X"12",X"49",X"92",X"A4",X"94",X"4A",X"2A",X"55",X"AA",X"52",X"55",X"A5",X"AA",
		X"5A",X"AD",X"AA",X"BA",X"54",X"4A",X"22",X"A4",X"A4",X"52",X"D5",X"AE",X"DF",X"B6",X"AD",X"55",
		X"AD",X"4A",X"55",X"55",X"55",X"55",X"A9",X"A4",X"2A",X"95",X"92",X"22",X"12",X"29",X"A5",X"94",
		X"AA",X"AA",X"AA",X"AA",X"14",X"49",X"94",X"92",X"AA",X"56",X"AB",X"55",X"55",X"AB",X"AA",X"52",
		X"2A",X"A9",X"A4",X"AA",X"AA",X"6A",X"55",X"55",X"2A",X"29",X"29",X"55",X"55",X"DD",X"D6",X"F6",
		X"ED",X"5A",X"A9",X"AA",X"AA",X"BE",X"DA",X"56",X"A9",X"94",X"54",X"55",X"55",X"55",X"95",X"48",
		X"A4",X"52",X"55",X"B5",X"56",X"55",X"55",X"95",X"AA",X"AA",X"B5",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"52",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"B5",
		X"AA",X"55",X"BF",X"6D",X"57",X"AB",X"9A",X"2A",X"95",X"4A",X"AA",X"52",X"A9",X"A4",X"28",X"29",
		X"49",X"4A",X"94",X"2A",X"55",X"55",X"55",X"55",X"B3",X"D6",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"52",X"55",X"55",X"55",X"55",X"55",X"55",X"AD",X"6A",X"55",X"AD",X"53",X"55",X"D5",X"DB",
		X"B6",X"6D",X"DB",X"BA",X"AD",X"AD",X"A5",X"4A",X"A9",X"52",X"95",X"A4",X"44",X"A5",X"14",X"89",
		X"94",X"24",X"A9",X"94",X"AA",X"AA",X"AA",X"56",X"AB",X"5A",X"55",X"AB",X"AA",X"AA",X"4A",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AD",X"AD",X"AA",X"AA",X"AA",X"AA",X"5A",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"95",X"54",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"D5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"4A",X"A5",X"4A",X"A9",X"AA",X"2A",X"C1",X"1D",X"E7",X"AD",X"D3",X"AE",X"76",X"55",
		X"EB",X"EA",X"5A",X"E6",X"38",X"82",X"6F",X"4F",X"39",X"8E",X"9A",X"31",X"CE",X"32",X"63",X"16",
		X"B3",X"91",X"09",X"73",X"E6",X"EB",X"62",X"E2",X"02",X"67",X"E7",X"1A",X"C7",X"E4",X"C8",X"CC",
		X"99",X"99",X"89",X"98",X"99",X"69",X"C4",X"98",X"29",X"87",X"99",X"33",X"E6",X"C4",X"CC",X"71",
		X"E6",X"CE",X"CC",X"39",X"C7",X"39",X"E7",X"EC",X"CC",X"98",X"E3",X"19",X"E3",X"26",X"C7",X"71",
		X"CC",X"66",X"8C",X"33",X"6F",X"CE",X"39",X"37",X"F3",X"6C",X"9E",X"79",X"8E",X"D9",X"8C",X"3B",
		X"8B",X"CC",X"18",X"8C",X"33",X"E3",X"0C",X"85",X"39",X"E6",X"0C",X"83",X"31",X"CE",X"4C",X"4C",
		X"1D",X"33",X"2E",X"1E",X"8F",X"39",X"E6",X"38",X"66",X"8E",X"9D",X"1C",X"33",X"37",X"66",X"1C",
		X"37",X"37",X"CE",X"0E",X"1E",X"C7",X"0E",X"3B",X"4E",X"2E",X"CE",X"C4",X"8D",X"1D",X"9A",X"19",
		X"26",X"CE",X"0D",X"66",X"CC",X"19",X"3D",X"E2",X"19",X"46",X"33",X"C7",X"1C",X"C5",X"71",X"8C",
		X"CB",X"11",X"9B",X"AC",X"46",X"4E",X"DC",X"B0",X"0E",X"66",X"C6",X"8C",X"EC",X"98",X"39",X"66",
		X"E5",X"89",X"99",X"1B",X"67",X"E6",X"C6",X"B8",X"C9",X"9D",X"F3",X"14",X"E7",X"1C",X"E7",X"8E",
		X"C7",X"1D",X"C7",X"35",X"9D",X"6A",X"C7",X"39",X"66",X"63",X"8C",X"93",X"59",X"66",X"C6",X"70",
		X"89",X"93",X"4E",X"47",X"C6",X"84",X"C7",X"5C",X"8C",X"E3",X"48",X"A3",X"2A",X"E7",X"30",X"C3",
		X"19",X"F5",X"D5",X"DA",X"C2",X"1B",X"37",X"F2",X"A1",X"5A",X"C3",X"CC",X"FA",X"A0",X"47",X"CE",
		X"D1",X"D0",X"CC",X"E1",X"21",X"35",X"E5",X"C8",X"58",X"71",X"51",X"35",X"EA",X"30",X"9D",X"72",
		X"EA",X"5C",X"F1",X"B2",X"5A",X"F1",X"C8",X"BC",X"B8",X"33",X"AE",X"D2",X"34",X"5C",X"E5",X"D4",
		X"9C",X"95",X"79",X"54",X"A5",X"4E",X"66",X"4E",X"F5",X"CA",X"1E",X"8A",X"AA",X"8D",X"AA",X"2A",
		X"5F",X"54",X"95",X"0E",X"C5",X"32",X"5A",X"52",X"55",X"AC",X"A4",X"55",X"AC",X"A2",X"2A",X"A1",
		X"A2",X"56",X"5A",X"4D",X"B5",X"4C",X"39",X"E5",X"EA",X"AE",X"D5",X"0E",X"D7",X"5A",X"55",X"27",
		X"5D",X"BA",X"56",X"BB",X"6E",X"AF",X"AA",X"A2",X"2A",X"AA",X"55",X"55",X"52",X"8A",X"AA",X"50",
		X"0D",X"55",X"92",X"2A",X"B5",X"94",X"AA",X"D4",X"95",X"AA",X"EA",X"AA",X"B4",X"88",X"EB",X"B0",
		X"52",X"AB",X"EA",X"A8",X"5A",X"A5",X"2A",X"BA",X"AA",X"54",X"54",X"54",X"A9",X"52",X"D5",X"B2",
		X"2A",X"AB",X"AA",X"45",X"D5",X"AA",X"A5",X"CA",X"25",X"5D",X"89",X"2E",X"6A",X"95",X"16",X"B5",
		X"2A",X"97",X"54",X"AD",X"16",X"57",X"55",X"59",X"1A",X"5F",X"AC",X"94",X"B6",X"BA",X"BA",X"BA",
		X"35",X"B5",X"92",X"7A",X"51",X"55",X"55",X"69",X"AA",X"D2",X"4A",X"51",X"55",X"A5",X"AA",X"AE",
		X"5E",X"52",X"55",X"AD",X"AA",X"7A",X"A9",X"8B",X"5E",X"A9",X"2B",X"AA",X"4A",X"2B",X"55",X"55",
		X"2B",X"55",X"8A",X"25",X"35",X"2A",X"A5",X"B4",X"4E",X"B5",X"5C",X"95",X"AA",X"A8",X"56",X"55",
		X"55",X"AD",X"D7",X"22",X"95",X"D2",X"5A",X"95",X"A4",X"AA",X"AA",X"AA",X"AA",X"AA",X"8B",X"5E",
		X"A9",X"55",X"AC",X"AA",X"56",X"55",X"55",X"55",X"15",X"AD",X"AA",X"0A",X"55",X"55",X"55",X"A5",
		X"AA",X"5A",X"45",X"55",X"AA",X"17",X"AD",X"AA",X"7A",X"5D",X"5B",X"6D",X"AB",X"5B",X"95",X"2E",
		X"59",X"55",X"95",X"54",X"49",X"95",X"2A",X"AA",X"A2",X"AA",X"AA",X"AA",X"AA",X"AA",X"56",X"E9",
		X"AA",X"D2",X"2A",X"D5",X"AA",X"D6",X"AA",X"A2",X"AA",X"4A",X"55",X"52",X"55",X"55",X"55",X"55",
		X"55",X"55",X"95",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"AF",X"54",X"8B",X"6A",X"A9",X"AA",
		X"AA",X"95",X"AA",X"AA",X"AA",X"A2",X"A2",X"AA",X"92",X"4A",X"55",X"D5",X"AA",X"B5",X"AA",X"AA",
		X"AA",X"AA",X"6A",X"A9",X"AA",X"5A",X"97",X"94",X"AA",X"AA",X"AA",X"8A",X"AA",X"52",X"55",X"29",
		X"55",X"15",X"AA",X"AA",X"56",X"55",X"AB",X"AE",X"55",X"7D",X"D5",X"3D",X"F4",X"8A",X"5B",X"A9",
		X"AA",X"AA",X"2A",X"55",X"55",X"55",X"AA",X"4A",X"55",X"55",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"56",X"D5",X"2A",X"5A",X"45",X"55",X"AA",X"AA",X"54",X"A5",X"AA",X"54",X"95",X"50",
		X"15",X"55",X"52",X"A9",X"AA",X"6A",X"AB",X"AA",X"AA",X"5A",X"55",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"55",X"AF",X"AA",X"55",X"55",X"55",X"55",X"55",X"AD",X"FA",
		X"55",X"77",X"B5",X"AD",X"6A",X"8B",X"AA",X"5F",X"55",X"55",X"55",X"55",X"95",X"4A",X"4A",X"A2",
		X"92",X"A4",X"4A",X"A9",X"AA",X"AA",X"75",X"55",X"75",X"55",X"55",X"55",X"AB",X"AA",X"92",X"AA",
		X"54",X"55",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"DA",X"AA",X"AA",X"AD",X"AA",X"AA",X"AA",
		X"4A",X"55",X"55",X"55",X"B5",X"AA",X"AA",X"AA",X"AA",X"4A",X"AA",X"A8",X"AA",X"54",X"25",X"AA",
		X"A4",X"AA",X"AA",X"AA",X"AA",X"AA",X"54",X"AB",X"AA",X"55",X"55",X"D5",X"AA",X"EA",X"95",X"AA",
		X"AA",X"AA",X"4A",X"55",X"55",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AE",X"AA",X"AA",X"AA",
		X"4A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"A5",X"AA",X"AA",X"AA",X"AA",X"55",X"75",X"55",X"AD",X"52",X"FB",X"52",X"55",X"AA",
		X"AA",X"56",X"55",X"55",X"D5",X"97",X"52",X"55",X"55",X"55",X"AA",X"AA",X"AA",X"DA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"4A",X"A9",X"AA",X"AA",X"AA",X"5A",X"55",X"55",X"54",X"15",X"AA",X"24",X"15",
		X"AA",X"4A",X"55",X"55",X"AB",X"5A",X"69",X"55",X"55",X"55",X"55",X"AB",X"AA",X"BA",X"AA",X"AA",
		X"2A",X"55",X"55",X"55",X"AB",X"AA",X"56",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"75",
		X"4B",X"55",X"55",X"55",X"55",X"55",X"55",X"A9",X"4A",X"55",X"52",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"AA",X"AA",X"AA",X"AB",X"AA",X"AA",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"AD",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"B5",X"AA",X"AA",X"AA",X"AA",X"AA",X"A4",X"52",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"DB",X"AA",X"AA",X"BA",X"AD",X"54",X"55",X"7B",X"BB",X"D6",X"9A",
		X"4A",X"A5",X"AA",X"54",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"55",X"D5",X"5D",X"55",X"95",X"5A",
		X"55",X"55",X"55",X"55",X"55",X"49",X"55",X"55",X"AB",X"54",X"95",X"AA",X"4A",X"2A",X"55",X"95",
		X"54",X"55",X"55",X"55",X"AB",X"55",X"55",X"B5",X"EA",X"D7",X"B6",X"AD",X"54",X"55",X"95",X"AA",
		X"AA",X"92",X"AA",X"AA",X"AA",X"45",X"55",X"AB",X"AA",X"AA",X"BA",X"AA",X"6A",X"55",X"AB",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"54",X"4A",X"55",X"45",X"2A",X"89",X"2A",X"25",X"AA",X"54",X"55",
		X"55",X"55",X"55",X"55",X"D5",X"AE",X"BA",X"AA",X"EA",X"6D",X"AB",X"6D",X"BB",X"6A",X"AA",X"AA",
		X"AA",X"54",X"55",X"55",X"A5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"AA",X"AA",X"52",X"92",X"54",X"55",X"55",
		X"55",X"B5",X"AA",X"AD",X"AA",X"EA",X"54",X"55",X"55",X"BD",X"6B",X"AB",X"AA",X"52",X"95",X"AA",
		X"4A",X"AA",X"AA",X"AA",X"92",X"54",X"55",X"55",X"D5",X"6A",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"92",X"44",X"22",X"12",X"49",X"52",X"92",X"4A",X"AA",
		X"AA",X"AA",X"AB",X"B6",X"AA",X"56",X"55",X"55",X"7D",X"DB",X"DA",X"B6",X"B6",X"95",X"AA",X"AA",
		X"AA",X"4A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"95",X"4A",X"A9",X"2A",X"A5",X"22",X"49",X"22",X"92",X"24",X"4A",X"29",X"A9",X"AA",X"AA",
		X"DA",X"D6",X"EA",X"DB",X"ED",X"EE",X"6E",X"BB",X"B6",X"AA",X"2A",X"A9",X"4A",X"A9",X"94",X"94",
		X"4A",X"55",X"75",X"AD",X"EA",X"5B",X"D7",X"5A",X"D7",X"AA",X"15",X"84",X"24",X"92",X"A4",X"44",
		X"22",X"89",X"54",X"AA",X"AA",X"AA",X"52",X"55",X"6B",X"6F",X"5B",X"DB",X"DA",X"B6",X"B7",X"BB",
		X"DD",X"B6",X"AD",X"D6",X"D6",X"AA",X"56",X"AA",X"52",X"2A",X"A5",X"28",X"91",X"28",X"91",X"92",
		X"24",X"89",X"24",X"49",X"22",X"A9",X"94",X"54",X"55",X"44",X"55",X"A9",X"76",X"BF",X"7B",X"7F",
		X"FF",X"FF",X"57",X"25",X"21",X"52",X"B6",X"A2",X"44",X"20",X"A0",X"2A",X"B5",X"AA",X"52",X"52",
		X"AA",X"6A",X"B7",X"56",X"95",X"52",X"DD",X"BD",X"BB",X"B7",X"D6",X"5A",X"5B",X"DB",X"D6",X"AA",
		X"AA",X"A8",X"AA",X"AA",X"AA",X"AA",X"24",X"A5",X"94",X"4A",X"24",X"4A",X"24",X"52",X"52",X"52",
		X"92",X"92",X"52",X"55",X"55",X"55",X"55",X"B5",X"BA",X"7A",X"DB",X"DA",X"7A",X"DB",X"6D",X"6D",
		X"55",X"6B",X"A5",X"AA",X"52",X"95",X"2A",X"95",X"AA",X"94",X"A4",X"48",X"54",X"2A",X"A5",X"AA",
		X"02",X"00",X"A0",X"52",X"FF",X"FF",X"F7",X"56",X"6D",X"77",X"B7",X"DF",X"FF",X"01",X"40",X"00",
		X"90",X"B6",X"40",X"8A",X"00",X"21",X"6B",X"AA",X"6D",X"15",X"A9",X"AA",X"BA",X"F7",X"DD",X"F6",
		X"D6",X"76",X"5B",X"AB",X"EE",X"DF",X"FF",X"77",X"2B",X"AD",X"EA",X"EE",X"6E",X"6B",X"DB",X"FF",
		X"01",X"40",X"00",X"80",X"B6",X"00",X"89",X"00",X"40",X"96",X"A4",X"AA",X"2A",X"A4",X"55",X"55",
		X"7B",X"B7",X"76",X"AB",X"A9",X"BA",X"FB",X"FF",X"DF",X"B5",X"AA",X"DA",X"FB",X"F7",X"6E",X"AB",
		X"DE",X"FF",X"01",X"14",X"00",X"C0",X"3D",X"20",X"85",X"00",X"40",X"15",X"51",X"D5",X"0A",X"51",
		X"55",X"2A",X"ED",X"AD",X"52",X"ED",X"EE",X"76",X"B7",X"55",X"ED",X"FF",X"7E",X"F7",X"5D",X"75",
		X"FF",X"FF",X"01",X"0E",X"00",X"C1",X"3D",X"88",X"85",X"00",X"80",X"25",X"52",X"DA",X"0A",X"A9",
		X"52",X"8A",X"6A",X"55",X"FF",X"AA",X"AA",X"56",X"F5",X"FF",X"7F",X"B7",X"5B",X"7D",X"FF",X"FF",
		X"0F",X"60",X"00",X"08",X"EE",X"83",X"18",X"14",X"00",X"A8",X"48",X"65",X"5B",X"00",X"55",X"AB",
		X"D0",X"5E",X"A5",X"DA",X"EF",X"DE",X"7F",X"B7",X"FD",X"7F",X"F7",X"FF",X"03",X"30",X"08",X"80",
		X"FF",X"40",X"8A",X"02",X"00",X"15",X"24",X"ED",X"16",X"52",X"05",X"44",X"F6",X"DE",X"7D",X"55",
		X"6D",X"FF",X"EF",X"FF",X"FF",X"01",X"28",X"00",X"C0",X"7F",X"90",X"15",X"01",X"00",X"0B",X"92",
		X"EA",X"8D",X"E8",X"14",X"08",X"BA",X"DB",X"FD",X"2B",X"E9",X"FD",X"FE",X"FF",X"FF",X"0F",X"00",
		X"01",X"00",X"FC",X"07",X"6A",X"20",X"00",X"20",X"40",X"EA",X"3D",X"A1",X"02",X"20",X"B2",X"77",
		X"6F",X"AB",X"AA",X"F4",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"FF",X"40",X"85",X"02",X"00",
		X"00",X"BA",X"EF",X"0F",X"00",X"01",X"24",X"FD",X"5F",X"6D",X"55",X"4A",X"FF",X"FF",X"FF",X"03",
		X"00",X"00",X"80",X"FF",X"01",X"15",X"05",X"00",X"F8",X"6E",X"FF",X"17",X"00",X"00",X"91",X"FE",
		X"7F",X"A5",X"5A",X"6D",X"FF",X"FF",X"01",X"80",X"A4",X"F6",X"FF",X"B5",X"FB",X"8B",X"F4",X"26",
		X"42",X"29",X"00",X"00",X"95",X"24",X"55",X"00",X"00",X"00",X"52",X"FF",X"AF",X"DA",X"FB",X"FF",
		X"7F",X"00",X"00",X"80",X"FE",X"FF",X"FF",X"2F",X"90",X"BF",X"52",X"BB",X"25",X"00",X"00",X"22",
		X"A9",X"0A",X"00",X"00",X"00",X"72",X"FF",X"AF",X"F6",X"FB",X"FF",X"01",X"10",X"00",X"00",X"FF",
		X"81",X"15",X"15",X"A1",X"FF",X"BF",X"52",X"2F",X"02",X"20",X"04",X"50",X"92",X"48",X"15",X"00",
		X"FB",X"FD",X"0F",X"00",X"FD",X"FF",X"C1",X"2F",X"00",X"00",X"54",X"F9",X"FF",X"4F",X"E8",X"3F",
		X"D2",X"FF",X"02",X"40",X"05",X"48",X"ED",X"22",X"AA",X"A4",X"DA",X"FF",X"FF",X"FF",X"3F",X"00",
		X"20",X"00",X"D8",X"97",X"D4",X"7F",X"05",X"F8",X"7F",X"E5",X"FF",X"01",X"AA",X"02",X"00",X"AE",
		X"00",X"5A",X"00",X"AA",X"75",X"B5",X"FF",X"55",X"ED",X"56",X"EA",X"FF",X"DD",X"EE",X"B6",X"4A",
		X"48",X"D5",X"AA",X"6E",X"15",X"48",X"5F",X"64",X"5F",X"1B",X"A0",X"4D",X"00",X"00",X"00",X"D8",
		X"EA",X"2A",X"42",X"00",X"EA",X"FF",X"BF",X"FF",X"1F",X"00",X"E0",X"B7",X"FF",X"3F",X"40",X"FF",
		X"AA",X"FF",X"3F",X"00",X"02",X"80",X"FD",X"7F",X"F5",X"1F",X"00",X"B5",X"26",X"F9",X"3F",X"F9",
		X"FF",X"07",X"00",X"00",X"E8",X"FF",X"FF",X"36",X"10",X"F5",X"FF",X"FF",X"DF",X"84",X"B4",X"45",
		X"FC",X"7F",X"A5",X"F7",X"02",X"F4",X"5F",X"F5",X"FF",X"A5",X"FE",X"3F",X"00",X"00",X"80",X"FE",
		X"BF",X"FF",X"13",X"FD",X"FF",X"FF",X"0B",X"00",X"00",X"A0",X"FF",X"6F",X"02",X"00",X"00",X"80",
		X"EA",X"FF",X"BB",X"DB",X"FF",X"07",X"E0",X"00",X"00",X"FF",X"E8",X"FF",X"01",X"E8",X"FB",X"FE",
		X"FF",X"17",X"28",X"00",X"60",X"BF",X"12",X"25",X"00",X"00",X"20",X"FA",X"FF",X"B6",X"ED",X"FF",
		X"07",X"E0",X"01",X"00",X"7E",X"00",X"FF",X"00",X"00",X"1B",X"FC",X"FF",X"EF",X"34",X"00",X"F0",
		X"A4",X"ED",X"1F",X"00",X"16",X"40",X"FF",X"FF",X"FF",X"07",X"00",X"00",X"00",X"DA",X"12",X"20",
		X"0B",X"00",X"FE",X"FF",X"DF",X"2F",X"00",X"08",X"82",X"FA",X"5B",X"55",X"09",X"20",X"FD",X"F7",
		X"FF",X"4F",X"2A",X"00",X"00",X"BD",X"EA",X"EF",X"24",X"00",X"A8",X"FF",X"FF",X"7F",X"55",X"01",
		X"20",X"00",X"40",X"AA",X"00",X"01",X"10",X"A1",X"FF",X"4F",X"94",X"00",X"F2",X"FF",X"FF",X"FF",
		X"0F",X"00",X"00",X"A0",X"FF",X"7F",X"B4",X"FF",X"51",X"FF",X"0B",X"00",X"01",X"00",X"B9",X"08",
		X"69",X"02",X"F4",X"5D",X"DB",X"FF",X"FF",X"03",X"A0",X"03",X"00",X"5D",X"00",X"FC",X"9F",X"F4",
		X"9F",X"F4",X"FF",X"D7",X"FF",X"06",X"70",X"01",X"00",X"48",X"20",X"2D",X"02",X"49",X"01",X"F0",
		X"5F",X"F5",X"FF",X"AF",X"FF",X"0F",X"00",X"00",X"00",X"FA",X"DA",X"BF",X"01",X"FC",X"FF",X"FE",
		X"FF",X"01",X"4C",X"00",X"80",X"24",X"20",X"4B",X"20",X"D2",X"4A",X"FA",X"FF",X"FF",X"FF",X"02",
		X"80",X"5B",X"A8",X"2E",X"01",X"68",X"AB",X"EE",X"FF",X"FF",X"FF",X"49",X"FF",X"02",X"AA",X"00",
		X"00",X"00",X"00",X"90",X"80",X"B4",X"0A",X"D9",X"3F",X"E0",X"7F",X"C0",X"FF",X"FF",X"03",X"00",
		X"00",X"E0",X"7F",X"FA",X"FF",X"00",X"FE",X"FF",X"FF",X"7F",X"80",X"05",X"00",X"00",X"00",X"80",
		X"08",X"00",X"A0",X"90",X"F7",X"5D",X"D2",X"DF",X"FE",X"FF",X"81",X"00",X"00",X"50",X"9B",X"F6",
		X"6E",X"55",X"BF",X"FF",X"FF",X"6F",X"F5",X"4E",X"88",X"94",X"00",X"00",X"00",X"00",X"00",X"80",
		X"E8",X"2F",X"29",X"21",X"11",X"EA",X"FE",X"FF",X"FF",X"07",X"00",X"F0",X"FE",X"FF",X"BF",X"FF",
		X"BF",X"EF",X"5F",X"A5",X"16",X"00",X"C0",X"0B",X"C8",X"02",X"00",X"00",X"00",X"E8",X"13",X"EC",
		X"4B",X"FA",X"FF",X"B7",X"FF",X"FF",X"FF",X"BF",X"50",X"D7",X"FD",X"FF",X"B7",X"FF",X"5B",X"FF",
		X"6F",X"ED",X"4F",X"00",X"00",X"00",X"50",X"05",X"B4",X"05",X"00",X"00",X"00",X"A0",X"11",X"D4",
		X"8A",X"F4",X"FF",X"FD",X"FF",X"FF",X"FF",X"BF",X"EA",X"FF",X"F6",X"FF",X"EF",X"DE",X"55",X"FF",
		X"BF",X"76",X"AB",X"4A",X"09",X"00",X"00",X"14",X"20",X"57",X"00",X"00",X"00",X"00",X"00",X"A2",
		X"AA",X"24",X"FD",X"FF",X"FD",X"FF",X"FF",X"55",X"D4",X"FE",X"FF",X"FF",X"FF",X"7D",X"DF",X"7B",
		X"FF",X"AD",X"B6",X"55",X"24",X"02",X"00",X"70",X"01",X"6A",X"01",X"A8",X"00",X"00",X"00",X"00",
		X"A8",X"44",X"6A",X"B7",X"EE",X"FF",X"FF",X"02",X"00",X"74",X"FF",X"FF",X"BF",X"FB",X"BB",X"FB",
		X"FF",X"77",X"B7",X"89",X"08",X"00",X"A8",X"AD",X"52",X"49",X"88",X"00",X"00",X"44",X"24",X"A2",
		X"54",X"22",X"FD",X"5F",X"FD",X"FF",X"01",X"48",X"80",X"FC",X"BF",X"EE",X"B7",X"A8",X"BF",X"FF",
		X"FF",X"6F",X"D5",X"AA",X"54",X"55",X"11",X"88",X"02",X"00",X"00",X"00",X"04",X"04",X"29",X"29",
		X"6A",X"77",X"FB",X"FF",X"87",X"20",X"08",X"A8",X"EF",X"5A",X"DB",X"25",X"20",X"F5",X"FF",X"FF",
		X"FF",X"FF",X"B7",X"AA",X"8A",X"A0",X"52",X"55",X"24",X"04",X"91",X"EE",X"ED",X"56",X"A9",X"EA",
		X"05",X"00",X"00",X"00",X"B4",X"80",X"28",X"49",X"50",X"D7",X"FA",X"FF",X"EF",X"FF",X"77",X"BB",
		X"26",X"92",X"48",X"AA",X"55",X"4A",X"6D",X"DB",X"77",X"DD",X"FF",X"09",X"FA",X"26",X"00",X"0A",
		X"00",X"50",X"5B",X"F5",X"37",X"C9",X"FE",X"6B",X"FF",X"57",X"7B",X"AF",X"B5",X"0A",X"40",X"09",
		X"00",X"29",X"00",X"A8",X"92",X"A4",X"56",X"55",X"55",X"15",X"52",X"57",X"4A",X"7F",X"B7",X"FD",
		X"EF",X"FE",X"BF",X"DF",X"B7",X"FD",X"B6",X"B6",X"2A",X"89",X"28",X"41",X"00",X"08",X"00",X"00",
		X"20",X"AD",X"92",X"A4",X"AA",X"AA",X"7F",X"B5",X"DD",X"6F",X"FB",X"DF",X"FB",X"7E",X"AB",X"05",
		X"00",X"A4",X"54",X"FB",X"56",X"5B",X"BB",X"EA",X"BF",X"00",X"48",X"15",X"A8",X"5D",X"81",X"54",
		X"01",X"20",X"09",X"54",X"5B",X"A5",X"FE",X"97",X"FA",X"BF",X"F6",X"FF",X"A0",X"FF",X"45",X"BB",
		X"0A",X"AA",X"25",X"80",X"56",X"00",X"52",X"08",X"6A",X"AB",X"A8",X"AF",X"92",X"EE",X"A5",X"EE",
		X"5B",X"65",X"57",X"A2",X"FF",X"03",X"6A",X"05",X"00",X"48",X"40",X"BD",X"55",X"D5",X"6D",X"ED",
		X"FF",X"BE",X"6D",X"77",X"DB",X"37",X"49",X"DD",X"45",X"54",X"01",X"A8",X"05",X"40",X"2A",X"40",
		X"AD",X"0A",X"69",X"0B",X"D9",X"2D",X"01",X"6D",X"05",X"A9",X"54",X"F5",X"77",X"FF",X"B5",X"7B",
		X"FF",X"BA",X"6F",X"B7",X"BD",X"B7",X"DA",X"AA",X"04",X"24",X"81",X"B4",X"15",X"29",X"05",X"00",
		X"00",X"00",X"2A",X"09",X"54",X"09",X"51",X"AD",X"DA",X"FF",X"FF",X"F6",X"6F",X"F7",X"BF",X"ED",
		X"B6",X"92",X"D4",X"4A",X"DD",X"4A",X"49",X"25",X"D2",X"4A",X"0A",X"20",X"00",X"21",X"22",X"90",
		X"2A",X"A9",X"44",X"A9",X"EE",X"6D",X"B7",X"7D",X"DF",X"DF",X"BE",X"AB",X"AA",X"12",X"6A",X"B7",
		X"56",X"D5",X"5A",X"89",X"FA",X"0A",X"91",X"08",X"00",X"22",X"92",X"22",X"A5",X"94",X"22",X"91",
		X"DA",X"FF",X"EB",X"AE",X"B6",X"FB",X"BF",X"F7",X"B6",X"92",X"B6",X"55",X"DD",X"55",X"EA",X"2A",
		X"D4",X"B7",X"00",X"12",X"00",X"48",X"89",X"A8",X"AA",X"44",X"55",X"20",X"AA",X"6D",X"EF",X"AF",
		X"75",X"FF",X"DA",X"7E",X"55",X"A5",X"55",X"B2",X"B7",X"AA",X"B6",X"52",X"7B",X"55",X"55",X"01",
		X"00",X"82",X"90",X"AA",X"24",X"55",X"22",X"AA",X"D6",X"AA",X"2A",X"11",X"55",X"D7",X"FF",X"FF",
		X"BB",X"6A",X"95",X"48",X"B5",X"DB",X"BD",X"55",X"12",X"55",X"A1",X"EE",X"2F",X"50",X"09",X"00",
		X"24",X"49",X"B5",X"44",X"A4",X"92",X"A4",X"D6",X"AA",X"EF",X"56",X"EB",X"B6",X"AA",X"AA",X"EA",
		X"FF",X"FF",X"BF",X"55",X"AD",X"4A",X"D5",X"D6",X"6A",X"55",X"11",X"55",X"EB",X"7F",X"05",X"20",
		X"00",X"20",X"55",X"49",X"15",X"01",X"91",X"44",X"AA",X"AD",X"6A",X"AD",X"AA",X"DA",X"EE",X"B6",
		X"BB",X"55",X"AB",X"AA",X"FD",X"FF",X"FF",X"5E",X"6B",X"5B",X"25",X"6A",X"5B",X"55",X"AB",X"22",
		X"7B",X"05",X"00",X"00",X"10",X"49",X"A2",X"94",X"84",X"10",X"22",X"4A",X"55",X"AD",X"D6",X"B5",
		X"B6",X"B6",X"EE",X"EE",X"7D",X"B7",X"AD",X"B5",X"B5",X"DA",X"EE",X"BB",X"DB",X"D6",X"AE",X"DD",
		X"6D",X"B5",X"AA",X"2A",X"A2",X"54",X"55",X"03",X"00",X"00",X"80",X"48",X"12",X"49",X"22",X"44",
		X"94",X"52",X"B5",X"D6",X"BA",X"D6",X"6A",X"DB",X"EE",X"FD",X"EE",X"76",X"B7",X"DB",X"6D",X"6B",
		X"AD",X"D5",X"DA",X"AE",X"56",X"EB",X"5A",X"75",X"55",X"94",X"AA",X"AA",X"AA",X"88",X"52",X"09",
		X"00",X"00",X"40",X"48",X"24",X"52",X"12",X"89",X"24",X"A5",X"AA",X"AA",X"B5",X"6E",X"DB",X"EE",
		X"76",X"77",X"77",X"77",X"BB",X"BB",X"DD",X"DD",X"B6",X"56",X"AD",X"55",X"6B",X"AD",X"55",X"49",
		X"95",X"92",X"24",X"12",X"41",X"94",X"84",X"48",X"12",X"89",X"10",X"84",X"24",X"22",X"49",X"4A",
		X"92",X"22",X"4A",X"A9",X"4A",X"55",X"55",X"55",X"AB",X"DB",X"BD",X"BB",X"7B",X"EF",X"EE",X"EE",
		X"7B",X"D7",X"EE",X"B6",X"76",X"AB",X"AA",X"B6",X"B5",X"0A",X"21",X"10",X"44",X"22",X"11",X"89",
		X"48",X"92",X"24",X"A5",X"AA",X"AA",X"56",X"D5",X"D5",X"6A",X"BB",X"DB",X"B6",X"DB",X"DA",X"76",
		X"ED",X"EE",X"DA",X"56",X"55",X"45",X"55",X"55",X"95",X"88",X"24",X"89",X"2A",X"49",X"11",X"12",
		X"51",X"95",X"52",X"22",X"A5",X"A4",X"52",X"95",X"AA",X"AA",X"AA",X"55",X"A5",X"DE",X"D5",X"56",
		X"55",X"A9",X"D4",X"56",X"FD",X"56",X"54",X"55",X"55",X"55",X"29",X"A9",X"5A",X"55",X"55",X"AA",
		X"DB",X"A5",X"EA",X"15",X"D5",X"2A",X"6A",X"5F",X"51",X"55",X"A9",X"5A",X"A5",X"2A",X"51",X"15",
		X"52",X"95",X"A8",X"AA",X"2A",X"A9",X"2A",X"54",X"55",X"55",X"AB",X"A4",X"AA",X"A8",X"5D",X"45",
		X"B5",X"AA",X"BF",X"55",X"75",X"AB",X"EE",X"55",X"A2",X"95",X"6A",X"5F",X"55",X"AA",X"90",X"AA",
		X"4A",X"75",X"41",X"6A",X"45",X"5A",X"95",X"54",X"25",X"AA",X"95",X"D4",X"5A",X"8A",X"AA",X"AA",
		X"54",X"2B",X"52",X"5D",X"45",X"FD",X"0A",X"ED",X"55",X"D4",X"A9",X"AA",X"57",X"95",X"BA",X"52",
		X"55",X"55",X"A5",X"2A",X"55",X"A9",X"AA",X"A5",X"AA",X"AA",X"52",X"D5",X"2A",X"B5",X"85",X"FA",
		X"15",X"BD",X"4A",X"56",X"A5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C5",
		X"4F",X"C6",X"00",X"F7",X"78",X"00",X"20",X"FB",X"86",X"01",X"20",X"F5",X"86",X"02",X"20",X"F1",
		X"FF",X"E8",X"FF",X"E8",X"FF",X"E8",X"FF",X"E0",X"FF",X"E8",X"FF",X"E8",X"FF",X"EC",X"FF",X"E8");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
