library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity joust2_bg_sound_bank_c is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of joust2_bg_sound_bank_c is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"B8",X"DD",X"19",X"0A",X"17",X"26",X"0A",X"96",X"16",X"97",X"17",X"0C",X"15",X"26",X"02",X"0C",
		X"14",X"12",X"86",X"14",X"B7",X"20",X"00",X"B6",X"40",X"00",X"C6",X"15",X"F7",X"20",X"01",X"DC",
		X"20",X"2B",X"1F",X"F7",X"60",X"00",X"54",X"4A",X"26",X"13",X"96",X"1F",X"B7",X"78",X"00",X"E6",
		X"A0",X"86",X"08",X"B7",X"78",X"00",X"10",X"9C",X"1D",X"25",X"02",X"86",X"FF",X"DD",X"20",X"F7",
		X"68",X"00",X"DC",X"19",X"3B",X"B6",X"5A",X"94",X"4A",X"95",X"AA",X"6D",X"AB",X"44",X"A4",X"A4",
		X"EA",X"DA",X"77",X"6B",X"55",X"83",X"88",X"92",X"52",X"D5",X"DA",X"7A",X"DB",X"56",X"B5",X"0A",
		X"A9",X"28",X"8A",X"AA",X"AA",X"AA",X"55",X"B5",X"BE",X"6D",X"75",X"55",X"15",X"25",X"45",X"8A",
		X"4A",X"A5",X"AA",X"5A",X"55",X"6F",X"B5",X"AE",X"AD",X"AA",X"AB",X"56",X"A2",X"AA",X"92",X"A2",
		X"A2",X"52",X"54",X"AA",X"54",X"55",X"55",X"AD",X"1E",X"AD",X"57",X"57",X"D5",X"56",X"2B",X"55",
		X"AA",X"4A",X"2A",X"55",X"C5",X"AA",X"A0",X"AA",X"AA",X"AA",X"AA",X"F4",X"4E",X"F5",X"55",X"85",
		X"AA",X"95",X"6A",X"BD",X"52",X"BC",X"C2",X"AA",X"AA",X"AA",X"C8",X"D2",X"AA",X"AA",X"6A",X"55",
		X"A4",X"AA",X"95",X"54",X"B5",X"6A",X"D5",X"AA",X"52",X"51",X"A9",X"7A",X"55",X"91",X"6A",X"55",
		X"55",X"17",X"1F",X"0A",X"BF",X"20",X"E9",X"57",X"11",X"AD",X"5E",X"55",X"52",X"55",X"95",X"AA",
		X"5E",X"28",X"7F",X"05",X"D5",X"2F",X"85",X"56",X"55",X"E5",X"55",X"A9",X"AB",X"AA",X"52",X"49",
		X"AB",X"54",X"AD",X"02",X"E9",X"AF",X"40",X"BA",X"5A",X"BC",X"56",X"D5",X"AA",X"AA",X"83",X"D2",
		X"AF",X"40",X"FC",X"15",X"A1",X"56",X"A5",X"5A",X"55",X"D5",X"7A",X"E1",X"BA",X"09",X"AA",X"BF",
		X"14",X"5A",X"75",X"2D",X"AA",X"45",X"F5",X"05",X"F8",X"2B",X"44",X"BE",X"0D",X"D0",X"BE",X"03",
		X"D5",X"17",X"D2",X"AE",X"81",X"DB",X"05",X"EA",X"5B",X"C0",X"7D",X"81",X"FA",X"52",X"72",X"D1",
		X"83",X"5B",X"07",X"56",X"BD",X"4A",X"89",X"D7",X"07",X"C9",X"DF",X"C0",X"FE",X"80",X"DA",X"56",
		X"49",X"74",X"2F",X"34",X"7D",X"50",X"7C",X"5D",X"D0",X"5E",X"60",X"79",X"AB",X"80",X"EE",X"0B",
		X"F8",X"0E",X"68",X"BD",X"AA",X"48",X"F5",X"03",X"AB",X"07",X"C5",X"BE",X"05",X"FC",X"0E",X"A8",
		X"3F",X"2C",X"1D",X"7A",X"0B",X"47",X"0F",X"47",X"AD",X"37",X"A0",X"FD",X"41",X"E8",X"0F",X"D4",
		X"2F",X"D0",X"AE",X"82",X"F6",X"0B",X"E8",X"1F",X"50",X"3F",X"50",X"ED",X"61",X"F1",X"A2",X"43",
		X"D7",X"06",X"56",X"37",X"F4",X"C0",X"55",X"07",X"8B",X"5F",X"05",X"FF",X"20",X"3D",X"A5",X"57",
		X"50",X"3F",X"19",X"DC",X"D6",X"C0",X"F2",X"87",X"F0",X"17",X"A8",X"6F",X"B0",X"BA",X"50",X"AB",
		X"07",X"EA",X"1B",X"A8",X"7E",X"41",X"7D",X"81",X"DA",X"0E",X"96",X"17",X"D1",X"0B",X"AF",X"40",
		X"BF",X"48",X"7D",X"81",X"FA",X"A2",X"BA",X"42",X"6B",X"E1",X"AE",X"20",X"EB",X"A5",X"BA",X"0A",
		X"3D",X"7A",X"1D",X"C8",X"F5",X"42",X"BD",X"82",X"53",X"FD",X"0A",X"5C",X"AF",X"42",X"DD",X"22",
		X"A1",X"7F",X"01",X"F6",X"07",X"EA",X"0B",X"78",X"AA",X"5E",X"C0",X"AF",X"50",X"BD",X"28",X"DC",
		X"05",X"E7",X"45",X"45",X"FB",X"0A",X"D8",X"3F",X"20",X"FD",X"02",X"D4",X"5F",X"E0",X"2F",X"48",
		X"FD",X"11",X"F2",X"1B",X"48",X"FF",X"02",X"FC",X"13",X"AA",X"97",X"05",X"FD",X"0B",X"B8",X"1E",
		X"C5",X"E8",X"FA",X"40",X"7D",X"A1",X"70",X"BD",X"05",X"EA",X"0F",X"C2",X"5F",X"10",X"FC",X"E2",
		X"70",X"E9",X"C0",X"5F",X"03",X"F6",X"61",X"D2",X"49",X"91",X"1F",X"1E",X"A3",X"1E",X"F4",X"AB",
		X"C0",X"AF",X"8A",X"1E",X"8B",X"7C",X"E1",X"53",X"F1",X"A0",X"3F",X"81",X"AF",X"49",X"4D",X"D1",
		X"FA",X"60",X"1E",X"A6",X"61",X"7B",X"01",X"F7",X"C1",X"1C",X"8A",X"3F",X"8C",X"47",X"3C",X"AC",
		X"27",X"A0",X"9F",X"C2",X"B3",X"08",X"FD",X"38",X"8E",X"E9",X"A0",X"FE",X"00",X"7F",X"19",X"BC",
		X"4A",X"F1",X"2B",X"E8",X"2F",X"81",X"FA",X"0F",X"D0",X"AF",X"50",X"DE",X"03",X"F4",X"1D",X"48",
		X"FF",X"00",X"7E",X"85",X"F1",X"2D",X"50",X"3F",X"41",X"FD",X"02",X"F4",X"17",X"D0",X"8F",X"0B",
		X"E8",X"C7",X"E1",X"0B",X"E8",X"07",X"EB",X"84",X"8F",X"73",X"0D",X"B4",X"1F",X"E0",X"73",X"1C",
		X"CE",X"07",X"F1",X"35",X"F4",X"85",X"E2",X"87",X"79",X"48",X"8F",X"EB",X"40",X"3F",X"8E",X"C1",
		X"7E",X"10",X"FE",X"80",X"F2",X"43",X"7C",X"8A",X"87",X"FC",X"30",X"3C",X"92",X"8F",X"3A",X"78",
		X"7C",X"01",X"FE",X"81",X"3E",X"E2",X"E1",X"7C",X"80",X"1F",X"8E",X"47",X"F2",X"1E",X"38",X"9F",
		X"22",X"BE",X"83",X"F3",X"70",X"3D",X"15",X"78",X"FC",X"00",X"3E",X"7C",X"81",X"9F",X"F0",X"03",
		X"F8",X"C3",X"78",X"0C",X"EF",X"C0",X"07",X"7E",X"A1",X"3B",X"E0",X"27",X"FC",X"0A",X"EC",X"03",
		X"B7",X"54",X"A3",X"7C",X"98",X"8E",X"AB",X"77",X"80",X"0F",X"6E",X"78",X"F8",X"38",X"F8",X"D0",
		X"0F",X"F0",X"E1",X"71",X"78",X"16",X"87",X"77",X"E0",X"AD",X"0E",X"EC",X"83",X"76",X"05",X"9F",
		X"40",X"DB",X"3E",X"40",X"1F",X"5E",X"C1",X"E3",X"F1",X"80",X"1F",X"3E",X"C0",X"0F",X"F5",X"01",
		X"7E",X"F0",X"03",X"F9",X"14",X"3E",X"C2",X"8F",X"C3",X"63",X"F8",X"03",X"3F",X"D0",X"27",X"FA",
		X"80",X"2F",X"3E",X"05",X"FD",X"C0",X"87",X"F8",X"92",X"1E",X"E4",X"F3",X"38",X"24",X"7F",X"80",
		X"4F",X"F0",X"71",X"0F",X"D4",X"87",X"0F",X"F0",X"83",X"C3",X"47",X"A9",X"0F",X"C5",X"F3",X"48",
		X"FE",X"01",X"FA",X"3C",X"04",X"3F",X"86",X"8F",X"E2",X"03",X"3F",X"84",X"1F",X"E3",X"E3",X"30",
		X"AE",X"0F",X"F0",X"13",X"BE",X"82",X"0F",X"F3",X"21",X"7C",X"0C",X"0F",X"C7",X"87",X"F1",X"11",
		X"3C",X"C6",X"C7",X"E0",X"33",X"3E",X"8E",X"E3",X"F8",X"40",X"FC",X"C0",X"AF",X"70",X"E8",X"3E",
		X"80",X"DF",X"C1",X"63",X"FA",X"30",X"3E",X"E0",X"C3",X"F8",X"18",X"3E",X"C6",X"C3",X"71",X"3C",
		X"3E",X"90",X"3F",X"F0",X"09",X"2F",X"1E",X"0F",X"D0",X"0F",X"F1",X"2B",X"1C",X"FA",X"41",X"F8",
		X"14",X"9E",X"87",X"96",X"1F",X"01",X"1F",X"5E",X"86",X"8F",X"CB",X"43",X"F4",X"63",X"78",X"18",
		X"8F",X"E3",X"41",X"3D",X"E5",X"47",X"3A",X"8E",X"0F",X"D0",X"07",X"3F",X"D4",X"C3",X"F1",X"01",
		X"1F",X"0F",X"0F",X"E5",X"03",X"3F",X"86",X"C7",X"E1",X"71",X"9C",X"F2",X"09",X"F8",X"44",X"1F",
		X"E2",X"61",X"3E",X"C4",X"C7",X"E3",X"C1",X"FA",X"C0",X"0F",X"F1",X"61",X"7C",X"98",X"E3",X"F8",
		X"82",X"FA",X"E0",X"C3",X"F0",X"38",X"1E",X"9C",X"C7",X"E1",X"C3",X"F0",X"C1",X"C7",X"E0",X"E3",
		X"78",X"1C",X"8E",X"BE",X"02",X"9E",X"FC",X"40",X"7C",X"F0",X"83",X"7C",X"3C",X"1E",X"5C",X"1E",
		X"3C",X"AC",X"07",X"FA",X"E0",X"78",X"F8",X"60",X"7C",X"78",X"09",X"3E",X"CF",X"03",X"FC",X"31",
		X"7C",X"28",X"1F",X"7C",X"38",X"1E",X"E3",X"C3",X"31",X"C7",X"43",X"D2",X"0F",X"1E",X"8E",X"07",
		X"1F",X"A3",X"C7",X"0F",X"E8",X"87",X"0F",X"8A",X"8F",X"23",X"A1",X"2F",X"7E",X"00",X"3F",X"3E",
		X"18",X"1E",X"87",X"63",X"55",X"F9",X"11",X"F8",X"EA",X"05",X"FD",X"88",X"0F",X"D4",X"7B",X"1C",
		X"A8",X"3F",X"18",X"1E",X"0F",X"CE",X"07",X"D5",X"8F",X"03",X"F9",X"83",X"7C",X"D0",X"C3",X"5D",
		X"A0",X"CF",X"87",X"C1",X"F3",X"E0",X"C3",X"E1",X"98",X"07",X"CE",X"0F",X"0F",X"D7",X"07",X"07",
		X"87",X"47",X"1D",X"38",X"8F",X"1E",X"C9",X"0F",X"0F",X"87",X"C7",X"15",X"1E",X"3E",X"5C",X"F4",
		X"1F",X"A0",X"7E",X"01",X"BC",X"0F",X"87",X"8F",X"83",X"87",X"C3",X"E3",X"88",X"A7",X"E1",X"C5",
		X"D0",X"E7",X"C1",X"F0",X"E1",X"E0",X"E3",X"F0",X"15",X"8C",X"1F",X"07",X"0F",X"0B",X"7E",X"1C",
		X"5E",X"0E",X"F8",X"79",X"38",X"3C",X"C2",X"CF",X"C1",X"C3",X"03",X"3F",X"0E",X"0F",X"2F",X"F8",
		X"71",X"78",X"78",X"E0",X"C7",X"C1",X"C3",X"0A",X"3F",X"0E",X"8F",X"53",X"F8",X"38",X"3C",X"2C",
		X"E1",X"C7",X"E1",X"F0",X"04",X"1F",X"87",X"C7",X"33",X"F8",X"38",X"3C",X"8E",X"E2",X"E3",X"70",
		X"38",X"87",X"8F",X"C3",X"E1",X"19",X"3E",X"07",X"8F",X"73",X"F8",X"38",X"3C",X"9C",X"E1",X"E3",
		X"F0",X"38",X"8E",X"8F",X"C3",X"E1",X"1C",X"1E",X"87",X"87",X"79",X"78",X"1C",X"1E",X"CE",X"F0",
		X"78",X"38",X"9C",X"C3",X"C3",X"E1",X"71",X"8C",X"8F",X"C3",X"E3",X"18",X"3E",X"0E",X"8F",X"63",
		X"3C",X"1C",X"1E",X"E3",X"F8",X"70",X"78",X"CC",X"E1",X"F1",X"F0",X"98",X"C3",X"C7",X"E1",X"71",
		X"8A",X"8F",X"C3",X"63",X"1C",X"1E",X"0F",X"87",X"1D",X"3C",X"1E",X"1E",X"F1",X"F0",X"70",X"78",
		X"6C",X"E1",X"F1",X"F0",X"88",X"87",X"87",X"C3",X"A3",X"07",X"8F",X"87",X"87",X"1E",X"1E",X"1E",
		X"1E",X"1F",X"3C",X"1C",X"3E",X"7C",X"F0",X"78",X"78",X"F8",X"E0",X"E1",X"E1",X"E1",X"83",X"87",
		X"C3",X"87",X"07",X"0F",X"C7",X"07",X"1F",X"1E",X"0E",X"3E",X"3C",X"3C",X"1C",X"3D",X"7C",X"78",
		X"38",X"7C",X"78",X"F0",X"70",X"F8",X"F0",X"C1",X"F1",X"D0",X"C3",X"83",X"C7",X"E1",X"C3",X"07",
		X"87",X"87",X"0F",X"0F",X"0F",X"8F",X"0F",X"2F",X"3C",X"1C",X"3E",X"3C",X"78",X"3C",X"3C",X"7C",
		X"F0",X"F0",X"F0",X"E1",X"C1",X"F1",X"D0",X"C3",X"83",X"C7",X"83",X"C7",X"07",X"8F",X"07",X"1F",
		X"1E",X"3C",X"1E",X"3C",X"3C",X"78",X"3C",X"F4",X"78",X"E0",X"F1",X"E0",X"E3",X"81",X"C7",X"C3",
		X"87",X"0B",X"1E",X"0F",X"3E",X"1E",X"3C",X"1E",X"7A",X"5C",X"F0",X"F1",X"E0",X"E1",X"C1",X"E3",
		X"A1",X"87",X"03",X"1F",X"0F",X"1E",X"0F",X"7C",X"1C",X"7A",X"B8",X"E0",X"E3",X"E1",X"C3",X"83",
		X"C7",X"61",X"87",X"0D",X"3E",X"1E",X"3E",X"3C",X"78",X"3C",X"7C",X"D8",X"E0",X"E3",X"C1",X"C7",
		X"83",X"C7",X"83",X"0F",X"17",X"7C",X"3C",X"78",X"3C",X"F0",X"74",X"F0",X"E1",X"81",X"C7",X"83",
		X"8F",X"07",X"1E",X"1E",X"3C",X"3E",X"F0",X"78",X"F0",X"E1",X"C1",X"C3",X"83",X"C7",X"07",X"3E",
		X"1E",X"3C",X"3C",X"F8",X"78",X"F0",X"F1",X"C0",X"C7",X"83",X"8F",X"07",X"1E",X"0F",X"3E",X"1E",
		X"78",X"3C",X"F8",X"F0",X"E0",X"C3",X"A1",X"C7",X"03",X"1F",X"0F",X"3E",X"3C",X"F0",X"78",X"F0",
		X"E1",X"81",X"8F",X"83",X"0F",X"0F",X"3E",X"1C",X"7C",X"78",X"F0",X"71",X"D0",X"E3",X"81",X"8F",
		X"07",X"1F",X"0F",X"3E",X"1C",X"FA",X"B8",X"E0",X"F1",X"E0",X"C3",X"83",X"8F",X"0B",X"1E",X"0F",
		X"7C",X"3C",X"F8",X"78",X"E0",X"E3",X"C1",X"87",X"07",X"3E",X"1E",X"3C",X"7A",X"E0",X"E3",X"E0",
		X"C3",X"05",X"1F",X"0F",X"3E",X"3C",X"78",X"3C",X"E8",X"E1",X"C1",X"C7",X"C1",X"0F",X"0F",X"1E",
		X"87",X"7A",X"3C",X"F8",X"78",X"F0",X"E1",X"C1",X"C7",X"41",X"1F",X"07",X"3E",X"1E",X"7C",X"78",
		X"F0",X"78",X"E0",X"C3",X"83",X"C7",X"83",X"1F",X"0E",X"3E",X"1C",X"FC",X"70",X"E0",X"E3",X"C1",
		X"87",X"07",X"0F",X"0F",X"3E",X"3C",X"78",X"3C",X"F8",X"F0",X"E0",X"C3",X"A1",X"0F",X"87",X"7C",
		X"0E",X"BE",X"78",X"F0",X"71",X"C8",X"C7",X"21",X"3E",X"87",X"3E",X"74",X"F8",X"38",X"E8",X"E3",
		X"C0",X"C7",X"E1",X"0B",X"0F",X"1E",X"1E",X"7A",X"78",X"F0",X"78",X"F8",X"C2",X"85",X"87",X"07",
		X"1F",X"1E",X"3C",X"1E",X"FA",X"F0",X"E0",X"F1",X"E0",X"87",X"03",X"8F",X"87",X"1E",X"1E",X"7C",
		X"3C",X"F8",X"F0",X"E0",X"E1",X"E1",X"C3",X"83",X"8F",X"07",X"1F",X"1E",X"78",X"3C",X"F8",X"F0",
		X"E0",X"E3",X"E0",X"87",X"03",X"8F",X"87",X"1E",X"1E",X"7C",X"1C",X"FC",X"70",X"F0",X"F1",X"E0",
		X"43",X"87",X"8F",X"83",X"1E",X"1E",X"3C",X"1E",X"7C",X"E8",X"F0",X"F1",X"E0",X"C3",X"83",X"C7",
		X"C3",X"87",X"1E",X"3E",X"0E",X"3E",X"78",X"F0",X"78",X"F8",X"A0",X"C3",X"E3",X"C1",X"07",X"0F",
		X"8F",X"C3",X"47",X"3C",X"3C",X"1E",X"3C",X"78",X"F8",X"38",X"7C",X"C8",X"E1",X"E3",X"E0",X"83",
		X"87",X"0F",X"87",X"0F",X"39",X"3E",X"1C",X"7C",X"E8",X"F0",X"38",X"F8",X"44",X"C7",X"C7",X"C1",
		X"47",X"0E",X"8F",X"83",X"CF",X"78",X"78",X"78",X"78",X"E8",X"E1",X"71",X"F8",X"18",X"0F",X"8F",
		X"83",X"47",X"0D",X"8F",X"83",X"C7",X"E2",X"F1",X"38",X"78",X"B4",X"F2",X"30",X"7C",X"0C",X"8F",
		X"87",X"C3",X"87",X"0D",X"8F",X"C3",X"C7",X"F0",X"78",X"1C",X"3C",X"AE",X"F8",X"18",X"7C",X"8C",
		X"C7",X"E3",X"E1",X"71",X"85",X"8F",X"83",X"C7",X"71",X"78",X"1C",X"1E",X"97",X"E8",X"38",X"78",
		X"1C",X"87",X"C7",X"E1",X"E1",X"14",X"8F",X"87",X"C7",X"71",X"78",X"1C",X"1E",X"1E",X"F1",X"78",
		X"78",X"1C",X"87",X"C7",X"C3",X"D1",X"25",X"8F",X"83",X"A7",X"69",X"78",X"1E",X"8E",X"2E",X"F1",
		X"38",X"BC",X"2A",X"83",X"E7",X"E1",X"F0",X"22",X"8F",X"C3",X"E3",X"38",X"78",X"0E",X"0F",X"8F",
		X"F0",X"1C",X"3C",X"8D",X"C3",X"E3",X"70",X"BC",X"0A",X"C7",X"E3",X"B1",X"38",X"3C",X"0F",X"87",
		X"57",X"70",X"1E",X"5E",X"CA",X"E1",X"71",X"38",X"3D",X"86",X"73",X"78",X"55",X"0C",X"9F",X"C3",
		X"D9",X"2A",X"1C",X"8F",X"57",X"E1",X"F0",X"38",X"8E",X"8B",X"83",X"D3",X"BC",X"03",X"0E",X"CF",
		X"61",X"5E",X"1C",X"9C",X"E3",X"2B",X"F0",X"F0",X"2C",X"C7",X"83",X"63",X"0E",X"5F",X"0B",X"0E",
		X"1F",X"E3",X"7A",X"F0",X"70",X"F8",X"5C",X"F0",X"F0",X"38",X"2E",X"0F",X"3E",X"06",X"EF",X"4A",
		X"28",X"9F",X"A1",X"DB",X"E0",X"F0",X"78",X"78",X"58",X"C1",X"E7",X"70",X"33",X"0E",X"1E",X"87",
		X"0F",X"19",X"7C",X"16",X"77",X"E1",X"E0",X"B3",X"78",X"11",X"87",X"8F",X"53",X"2F",X"1C",X"3C",
		X"87",X"2F",X"E1",X"F0",X"69",X"EC",X"0A",X"C3",X"33",X"FA",X"14",X"1C",X"3E",X"C7",X"D5",X"70",
		X"AC",X"E1",X"D7",X"C0",X"C3",X"E3",X"70",X"3C",X"1C",X"1E",X"7C",X"17",X"78",X"F8",X"0C",X"1E",
		X"87",X"87",X"93",X"F5",X"0C",X"3C",X"3E",X"96",X"4B",X"38",X"3C",X"1E",X"3E",X"A3",X"D4",X"33",
		X"7C",X"2A",X"1C",X"9E",X"C3",X"A7",X"30",X"3E",X"83",X"6F",X"A1",X"E2",X"33",X"F8",X"18",X"1E",
		X"8F",X"C3",X"57",X"38",X"9C",X"43",X"AF",X"E0",X"E2",X"31",X"7C",X"16",X"C6",X"33",X"F9",X"0A",
		X"3C",X"3C",X"07",X"CF",X"C1",X"99",X"C3",X"D7",X"82",X"C3",X"E7",X"F0",X"38",X"1A",X"CF",X"E2",
		X"2B",X"78",X"F8",X"1C",X"1E",X"87",X"C3",X"E3",X"F8",X"10",X"0F",X"8F",X"C3",X"E3",X"38",X"1C",
		X"C7",X"97",X"E0",X"E1",X"39",X"3C",X"1C",X"17",X"4E",X"3E",X"07",X"1E",X"1E",X"87",X"8F",X"83",
		X"C7",X"E1",X"BA",X"14",X"7C",X"1C",X"3E",X"1C",X"1E",X"0F",X"8F",X"87",X"86",X"8F",X"C3",X"73",
		X"2C",X"9C",X"46",X"5F",X"61",X"8F",X"87",X"E3",X"A1",X"78",X"34",X"7A",X"2E",X"78",X"78",X"1C",
		X"1E",X"2E",X"7C",X"0C",X"CF",X"C3",X"E1",X"71",X"F8",X"18",X"1E",X"1E",X"96",X"47",X"93",X"1E",
		X"87",X"C7",X"61",X"F1",X"38",X"7C",X"94",X"87",X"C7",X"F1",X"51",X"1C",X"8F",X"C3",X"E3",X"70",
		X"78",X"1C",X"3E",X"C5",X"C3",X"39",X"7C",X"0C",X"0F",X"8F",X"C3",X"73",X"38",X"1E",X"87",X"C7",
		X"E1",X"F0",X"38",X"3C",X"8E",X"C3",X"71",X"78",X"0E",X"1E",X"1E",X"87",X"C7",X"78",X"38",X"8D",
		X"C7",X"C1",X"C3",X"79",X"78",X"1C",X"87",X"D3",X"F8",X"2C",X"3C",X"3C",X"0E",X"CF",X"E1",X"78",
		X"0C",X"9F",X"83",X"87",X"67",X"F1",X"38",X"0E",X"C7",X"E2",X"39",X"78",X"38",X"87",X"8F",X"E1",
		X"71",X"0C",X"1F",X"87",X"87",X"47",X"F9",X"18",X"0E",X"CF",X"F0",X"71",X"38",X"3C",X"CA",X"8F",
		X"E1",X"78",X"14",X"9F",X"C1",X"8B",X"A3",X"7E",X"0C",X"8F",X"63",X"F8",X"0C",X"9E",X"1C",X"D5",
		X"C7",X"70",X"3C",X"8A",X"CF",X"E0",X"95",X"51",X"3F",X"A4",X"C6",X"51",X"7C",X"06",X"A7",X"43",
		X"F9",X"11",X"BA",X"19",X"EC",X"87",X"F0",X"C3",X"E1",X"3C",X"C6",X"E3",X"30",X"1E",X"87",X"CB",
		X"51",X"F9",X"0C",X"D6",X"0B",X"FA",X"19",X"EC",X"E1",X"38",X"1E",X"47",X"7A",X"C4",X"C7",X"51",
		X"EA",X"91",X"FA",X"14",X"F4",X"31",X"7C",X"0E",X"53",X"F8",X"88",X"C7",X"C3",X"38",X"96",X"D7",
		X"04",X"AD",X"0F",X"7A",X"3C",X"94",X"2F",X"D0",X"37",X"18",X"F7",X"A0",X"AE",X"47",X"D1",X"29",
		X"AF",X"03",X"E5",X"0F",X"E4",X"3B",X"28",X"BF",X"A0",X"6F",X"B0",X"F8",X"03",X"B9",X"87",X"C3",
		X"B3",X"AC",X"17",X"24",X"3F",X"A4",X"F5",X"84",X"F4",X"91",X"7C",X"03",X"2E",X"1F",X"D8",X"2E",
		X"2C",X"7E",X"A2",X"E3",X"38",X"F8",X"94",X"EB",X"41",X"C8",X"8F",X"94",X"9F",X"82",X"FA",X"21",
		X"DD",X"25",X"E8",X"0F",X"A9",X"AF",X"40",X"7D",X"45",X"F9",X"0C",X"B4",X"27",X"75",X"A7",X"40",
		X"BF",X"50",X"7D",X"05",X"F4",X"13",X"D5",X"27",X"50",X"3F",X"A4",X"BD",X"02",X"FA",X"45",X"D6",
		X"13",X"B0",X"3F",X"52",X"AF",X"02",X"ED",X"93",X"EA",X"15",X"D0",X"1F",X"2A",X"5F",X"81",X"FA",
		X"89",X"FA",X"12",X"E8",X"4F",X"64",X"AF",X"40",X"FD",X"48",X"7D",X"05",X"74",X"2F",X"D2",X"57",
		X"A0",X"F6",X"42",X"7D",X"05",X"B4",X"2F",X"54",X"AF",X"40",X"FD",X"88",X"7A",X"03",X"E9",X"1E",
		X"D2",X"37",X"90",X"EE",X"A1",X"FA",X"12",X"68",X"9F",X"A4",X"BB",X"40",X"EE",X"43",X"EA",X"0B",
		X"A4",X"3F",X"A4",X"BE",X"40",X"F6",X"43",X"DA",X"17",X"C8",X"7D",X"48",X"F7",X"02",X"B5",X"0F",
		X"E9",X"1D",X"90",X"FB",X"20",X"ED",X"05",X"6A",X"1F",X"A4",X"BD",X"40",X"F5",X"0B",X"F2",X"2D",
		X"A8",X"F6",X"10",X"DF",X"82",X"B2",X"37",X"A4",X"77",X"90",X"BA",X"87",X"F2",X"2E",X"48",X"D7",
		X"45",X"DE",X"0A",X"B1",X"79",X"98",X"DB",X"10",X"B5",X"1E",X"E5",X"35",X"14",X"AD",X"8F",X"74",
		X"1D",X"84",X"F6",X"43",X"5A",X"87",X"D0",X"FA",X"50",X"EE",X"22",X"54",X"3F",X"8A",X"F5",X"04",
		X"DA",X"1F",X"A2",X"3D",X"09",X"ED",X"87",X"D4",X"17",X"C1",X"ED",X"83",X"EC",X"0B",X"E1",X"7E",
		X"44",X"DE",X"22",X"74",X"3D",X"A2",X"EE",X"10",X"DA",X"2F",X"A4",X"37",X"82",X"EE",X"07",X"E9",
		X"2D",X"84",X"BB",X"83",X"F4",X"15",X"E2",X"B6",X"21",X"F5",X"06",X"69",X"F5",X"C2",X"3C",X"0B",
		X"E9",X"DA",X"A1",X"BC",X"06",X"E5",X"BC",X"61",X"3C",X"8E",X"74",X"B5",X"C6",X"72",X"8C",X"6A",
		X"39",X"8F",X"71",X"1C",X"53",X"59",X"BB",X"A2",X"78",X"8E",X"70",X"BD",X"84",X"D5",X"45",X"51",
		X"DB",X"83",X"4A",X"6F",X"41",X"BA",X"97",X"90",X"FA",X"0A",X"A4",X"BF",X"40",X"EB",X"78",X"1A",
		X"E4",X"B7",X"A0",X"BE",X"22",X"AD",X"A4",X"DE",X"44",X"DD",X"C2",X"BC",X"28",X"BD",X"2A",X"B6",
		X"8A",X"E5",X"B2",X"54",X"A5",X"BA",X"0A",X"D5",X"43",X"EE",X"82",X"FC",X"15",X"D4",X"AE",X"50",
		X"55",X"A9",X"96",X"86",X"65",X"3D",X"A2",X"DA",X"2B",X"A4",X"57",X"A1",X"6A",X"55",X"95",X"AA",
		X"55",X"25",X"B5",X"AA",X"54",X"7D",X"2D",X"2A",X"5F",X"0B",X"D5",X"AD",X"90",X"B5",X"AB",X"A4",
		X"3A",X"25",X"55",X"AB",X"52",X"55",X"AA",X"56",X"85",X"D6",X"A2",X"6A",X"55",X"A8",X"AA",X"AA",
		X"2A",X"95",X"AA",X"56",X"A9",X"AB",X"50",X"75",X"15",X"55",X"2B",X"B5",X"4A",X"A9",X"AB",X"A8",
		X"BA",X"AA",X"68",X"AD",X"AB",X"B6",X"55",X"AA",X"4A",X"55",X"AB",X"8A",X"AA",X"AB",X"4A",X"55",
		X"55",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"25",X"AA",X"AA",X"AA",X"54",X"95",X"AA",X"55",X"55",
		X"D5",X"0B",X"A9",X"AE",X"2A",X"AD",X"4A",X"55",X"A5",X"AA",X"AA",X"AA",X"D5",X"AA",X"AA",X"BA",
		X"52",X"5B",X"15",X"AD",X"56",X"A5",X"AA",X"B8",X"AA",X"54",X"AA",X"56",X"55",X"55",X"25",X"51",
		X"EB",X"52",X"B5",X"A8",X"B4",X"AA",X"AA",X"AA",X"2A",X"2D",X"55",X"55",X"54",X"AB",X"2A",X"5D",
		X"D1",X"B4",X"AA",X"D6",X"A9",X"E8",X"AA",X"54",X"AA",X"AA",X"AA",X"AA",X"AA",X"D2",X"BA",X"6A",
		X"55",X"95",X"AA",X"AE",X"AA",X"2A",X"A9",X"6A",X"55",X"55",X"25",X"5A",X"BF",X"52",X"AA",X"AA",
		X"A4",X"AD",X"2A",X"6A",X"55",X"51",X"55",X"A9",X"AA",X"AB",X"4A",X"A5",X"D5",X"AA",X"2A",X"A5",
		X"55",X"D5",X"A8",X"54",X"B5",X"BA",X"AA",X"50",X"75",X"55",X"55",X"25",X"52",X"57",X"55",X"4F",
		X"45",X"7B",X"B5",X"74",X"AD",X"74",X"AD",X"54",X"55",X"A9",X"AA",X"AA",X"A5",X"52",X"D5",X"AA",
		X"AA",X"54",X"AA",X"AA",X"AA",X"D2",X"A8",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"AA",X"AA",X"6A",
		X"B5",X"A8",X"AA",X"4A",X"55",X"B5",X"D2",X"EA",X"52",X"B5",X"AA",X"54",X"BB",X"8A",X"AA",X"AA",
		X"AA",X"55",X"55",X"A5",X"EA",X"EA",X"DB",X"2A",X"AA",X"AA",X"AA",X"AA",X"50",X"55",X"55",X"55",
		X"0B",X"AA",X"AA",X"54",X"15",X"4A",X"A7",X"A2",X"5A",X"15",X"5A",X"AB",X"52",X"55",X"AD",X"9E",
		X"AA",X"4A",X"A5",X"6A",X"55",X"A9",X"56",X"55",X"15",X"AD",X"AB",X"52",X"FB",X"2A",X"EA",X"B5",
		X"52",X"5D",X"55",X"B7",X"8A",X"AA",X"16",X"AD",X"96",X"8A",X"AA",X"AA",X"AA",X"56",X"A5",X"52",
		X"28",X"55",X"14",X"AD",X"8A",X"52",X"AB",X"D2",X"D5",X"A3",X"AA",X"4A",X"55",X"AB",X"AA",X"AA",
		X"54",X"55",X"D5",X"AA",X"56",X"55",X"55",X"55",X"55",X"4D",X"4B",X"55",X"AA",X"AB",X"AA",X"4A",
		X"55",X"AD",X"46",X"69",X"55",X"3D",X"AA",X"8A",X"56",X"4B",X"45",X"D5",X"52",X"55",X"55",X"A9",
		X"6A",X"29",X"A9",X"AD",X"A8",X"52",X"B5",X"AA",X"AA",X"A8",X"56",X"B7",X"AA",X"50",X"FB",X"55",
		X"A8",X"5A",X"55",X"5A",X"55",X"B9",X"7A",X"0E",X"8D",X"5E",X"4A",X"AB",X"2A",X"55",X"AD",X"4A",
		X"AB",X"0B",X"AF",X"4A",X"D7",X"56",X"51",X"55",X"95",X"AA",X"AA",X"54",X"55",X"AA",X"AA",X"A5",
		X"4A",X"D5",X"52",X"49",X"AA",X"6A",X"55",X"AA",X"36",X"AA",X"AE",X"96",X"AA",X"6A",X"B4",X"74",
		X"15",X"AA",X"AB",X"52",X"55",X"4B",X"D5",X"AA",X"6A",X"A9",X"AA",X"A7",X"AA",X"53",X"A9",X"1E",
		X"55",X"AD",X"AA",X"2A",X"5A",X"BA",X"54",X"5A",X"15",X"55",X"55",X"95",X"96",X"C2",X"52",X"45",
		X"75",X"2A",X"AA",X"56",X"07",X"FC",X"08",X"7F",X"C4",X"87",X"E3",X"03",X"7C",X"38",X"3E",X"8C",
		X"87",X"87",X"FE",X"C0",X"C3",X"F0",X"01",X"3F",X"D4",X"07",X"F8",X"61",X"3D",X"E0",X"C7",X"F0",
		X"23",X"7C",X"1C",X"1F",X"E1",X"C3",X"F8",X"21",X"1E",X"1C",X"0F",X"0F",X"0F",X"C7",X"E7",X"E0",
		X"E1",X"F8",X"80",X"3F",X"D4",X"03",X"7E",X"C8",X"1F",X"E2",X"43",X"F8",X"11",X"3E",X"9C",X"0F",
		X"E1",X"C3",X"F1",X"70",X"78",X"3C",X"CC",X"07",X"0F",X"C7",X"07",X"FC",X"21",X"3E",X"E2",X"83",
		X"F7",X"10",X"1F",X"C1",X"0F",X"F8",X"70",X"FC",X"08",X"0F",X"C7",X"87",X"F1",X"F0",X"78",X"3C",
		X"78",X"38",X"7E",X"80",X"0F",X"E3",X"07",X"DE",X"70",X"0F",X"F1",X"21",X"FD",X"80",X"1F",X"C3",
		X"C7",X"F8",X"70",X"7C",X"88",X"0F",X"C3",X"8F",X"F0",X"78",X"78",X"38",X"3C",X"1C",X"3F",X"E0",
		X"8F",X"F0",X"11",X"3F",X"D4",X"0F",X"F8",X"50",X"7E",X"88",X"8F",X"E3",X"43",X"7C",X"38",X"3E",
		X"C4",X"87",X"E3",X"43",X"3C",X"38",X"7C",X"84",X"87",X"C7",X"47",X"F8",X"70",X"7C",X"C0",X"0F",
		X"F5",X"03",X"7E",X"B0",X"0F",X"F1",X"E1",X"F8",X"80",X"1F",X"8E",X"8F",X"F8",X"70",X"7C",X"80",
		X"0F",X"C7",X"47",X"F8",X"30",X"7E",X"C0",X"0F",X"F9",X"23",X"7C",X"C8",X"1F",X"F0",X"43",X"F8",
		X"11",X"3F",X"8C",X"0F",X"F8",X"61",X"FC",X"80",X"0F",X"C7",X"47",X"FC",X"20",X"3F",X"E0",X"C7",
		X"F0",X"21",X"7E",X"C8",X"0F",X"F1",X"61",X"FC",X"88",X"0F",X"E1",X"47",X"FC",X"30",X"3E",X"E0",
		X"87",X"F8",X"11",X"3E",X"98",X"0F",X"F1",X"61",X"7C",X"88",X"1F",X"E2",X"07",X"FC",X"30",X"3E",
		X"C4",X"0F",X"FA",X"21",X"7C",X"14",X"3F",X"E2",X"07",X"FC",X"01",X"3E",X"8E",X"1F",X"E1",X"C3",
		X"F8",X"88",X"1F",X"D4",X"C7",X"F8",X"A0",X"3E",X"C4",X"0F",X"F1",X"23",X"7E",X"90",X"1F",X"E2",
		X"C3",X"F8",X"10",X"3F",X"E8",X"87",X"F8",X"41",X"3F",X"C4",X"0F",X"F2",X"43",X"7C",X"18",X"3F",
		X"C2",X"07",X"F5",X"21",X"3E",X"8C",X"0F",X"F1",X"83",X"7E",X"08",X"1F",X"E6",X"C7",X"F0",X"41",
		X"7E",X"88",X"1F",X"E2",X"47",X"F8",X"81",X"3F",X"C4",X"07",X"F3",X"23",X"7C",X"18",X"1F",X"C2",
		X"87",X"F9",X"21",X"3E",X"A8",X"0F",X"F1",X"83",X"7D",X"10",X"1F",X"DC",X"87",X"F8",X"41",X"3F",
		X"88",X"0F",X"EE",X"43",X"FC",X"E0",X"1F",X"E0",X"07",X"F7",X"10",X"3F",X"F8",X"83",X"F8",X"C1",
		X"0F",X"C6",X"0F",X"5E",X"3C",X"7C",X"C0",X"8F",X"C3",X"07",X"F9",X"21",X"7E",X"D0",X"0F",X"E1",
		X"83",X"FD",X"10",X"1F",X"AC",X"87",X"F8",X"C1",X"3D",X"C4",X"0F",X"7E",X"30",X"EE",X"78",X"E0",
		X"F0",X"F0",X"C1",X"E3",X"E1",X"83",X"87",X"F3",X"C1",X"07",X"3F",X"F0",X"83",X"1F",X"7C",X"F0",
		X"C1",X"0E",X"FC",X"81",X"0F",X"7E",X"E0",X"C1",X"0F",X"3E",X"F0",X"83",X"0F",X"7E",X"F0",X"83",
		X"1F",X"7C",X"E0",X"83",X"EB",X"F0",X"F0",X"11",X"F8",X"F0",X"A3",X"F0",X"E1",X"0B",X"E3",X"C2",
		X"87",X"0F",X"7E",X"E0",X"0F",X"3E",X"F8",X"81",X"1F",X"F8",X"C0",X"87",X"F5",X"E0",X"E1",X"07",
		X"F0",X"C3",X"3F",X"C0",X"07",X"EF",X"30",X"F6",X"F0",X"C1",X"71",X"E1",X"C1",X"C3",X"1F",X"F0",
		X"83",X"0F",X"DE",X"80",X"CF",X"85",X"E3",X"03",X"3F",X"84",X"0F",X"0F",X"1F",X"FC",X"A0",X"8F",
		X"C1",X"07",X"DF",X"10",X"3F",X"F8",X"C1",X"F0",X"83",X"2F",X"0C",X"1F",X"FC",X"E0",X"C3",X"03",
		X"FF",X"20",X"FC",X"60",X"3E",X"E0",X"C3",X"3B",X"C8",X"1B",X"1E",X"7C",X"F0",X"03",X"3F",X"F8",
		X"E0",X"0F",X"7E",X"E0",X"83",X"0F",X"F8",X"E0",X"83",X"8F",X"83",X"0F",X"7E",X"10",X"3E",X"38",
		X"FF",X"C0",X"87",X"CB",X"0E",X"3E",X"F0",X"07",X"F8",X"C1",X"0F",X"8E",X"0B",X"1F",X"3C",X"1C",
		X"3F",X"F0",X"F0",X"C1",X"07",X"87",X"07",X"FE",X"01",X"DE",X"38",X"0F",X"F0",X"C3",X"1F",X"4C",
		X"FA",X"03",X"1F",X"7E",X"F0",X"07",X"1F",X"FC",X"C0",X"0F",X"3E",X"F0",X"A1",X"FC",X"E0",X"F0",
		X"61",X"F0",X"17",X"F0",X"E1",X"07",X"FE",X"E0",X"07",X"3E",X"F8",X"81",X"0F",X"1F",X"D4",X"07",
		X"3E",X"FC",X"C0",X"0F",X"3E",X"F8",X"81",X"0F",X"3F",X"F0",X"C3",X"1F",X"FC",X"F0",X"07",X"3F",
		X"FC",X"C0",X"0F",X"3F",X"F8",X"C3",X"1B",X"F6",X"F0",X"83",X"3D",X"F8",X"C1",X"1F",X"7E",X"F0",
		X"87",X"0F",X"FC",X"E1",X"05",X"7F",X"78",X"C2",X"1F",X"BC",X"E1",X"0F",X"7E",X"F0",X"07",X"7F",
		X"F0",X"C1",X"1F",X"7C",X"F0",X"83",X"1F",X"FC",X"C0",X"07",X"3F",X"F0",X"C1",X"0F",X"7C",X"F0",
		X"03",X"1F",X"7E",X"E0",X"87",X"1F",X"F8",X"F0",X"03",X"3F",X"FC",X"E0",X"07",X"3F",X"F8",X"E1",
		X"07",X"7F",X"F8",X"C0",X"0F",X"7E",X"F0",X"C3",X"07",X"7E",X"F0",X"83",X"1F",X"3E",X"F0",X"83",
		X"1F",X"EE",X"F0",X"83",X"1F",X"7C",X"F0",X"87",X"0F",X"FE",X"F0",X"81",X"1F",X"FC",X"F0",X"87",
		X"0F",X"FC",X"E0",X"07",X"3F",X"7C",X"E0",X"0F",X"1F",X"FC",X"E1",X"03",X"3F",X"F8",X"E0",X"07",
		X"1F",X"F8",X"C1",X"07",X"3F",X"F8",X"81",X"0F",X"3F",X"F0",X"C1",X"0F",X"7E",X"F8",X"C1",X"0F",
		X"3E",X"F0",X"C3",X"07",X"7E",X"F8",X"C0",X"0F",X"7E",X"F0",X"C3",X"07",X"7E",X"F0",X"C1",X"1F",
		X"3E",X"F0",X"83",X"0F",X"FE",X"F0",X"83",X"1F",X"FC",X"E0",X"07",X"1F",X"FC",X"E1",X"07",X"3F",
		X"F8",X"E0",X"0F",X"1F",X"F8",X"E1",X"07",X"3E",X"F8",X"C0",X"0F",X"1F",X"F8",X"C1",X"07",X"7F",
		X"F8",X"C0",X"0F",X"3E",X"F0",X"83",X"0F",X"FC",X"E0",X"03",X"3F",X"F8",X"C0",X"0F",X"1F",X"F0",
		X"C1",X"0F",X"7C",X"F8",X"81",X"0F",X"3E",X"F0",X"C3",X"0F",X"7C",X"F8",X"81",X"0F",X"7E",X"F0",
		X"C3",X"07",X"FE",X"F0",X"81",X"1F",X"FC",X"E0",X"87",X"0F",X"FC",X"E0",X"07",X"3F",X"BC",X"E0",
		X"07",X"1F",X"FC",X"E1",X"05",X"7F",X"78",X"C1",X"0F",X"7E",X"F0",X"83",X"0F",X"FC",X"E0",X"03",
		X"1F",X"3C",X"1C",X"07",X"3F",X"F0",X"E1",X"07",X"3E",X"F8",X"81",X"07",X"3F",X"F0",X"E0",X"07",
		X"3E",X"FC",X"C0",X"07",X"3F",X"F8",X"E0",X"07",X"3F",X"FC",X"C0",X"07",X"3F",X"F8",X"E1",X"03",
		X"3F",X"F8",X"E0",X"0F",X"1F",X"F8",X"C3",X"0B",X"7E",X"F8",X"C0",X"0F",X"7E",X"F0",X"C3",X"07",
		X"7E",X"F8",X"C0",X"0F",X"3E",X"F0",X"83",X"0F",X"FC",X"F0",X"03",X"1F",X"7C",X"E0",X"83",X"0F",
		X"7C",X"F0",X"D0",X"1C",X"FC",X"C0",X"87",X"1F",X"F8",X"F0",X"03",X"1F",X"7E",X"E0",X"83",X"1F",
		X"FC",X"F0",X"83",X"1F",X"FC",X"E0",X"87",X"1F",X"FC",X"E0",X"83",X"3F",X"7C",X"E0",X"07",X"1F",
		X"FC",X"E1",X"05",X"3F",X"FC",X"E0",X"0F",X"2F",X"F8",X"E1",X"07",X"3E",X"F8",X"C1",X"0F",X"3F",
		X"F0",X"C1",X"0F",X"7E",X"F8",X"80",X"0F",X"5E",X"F0",X"83",X"0F",X"7C",X"F0",X"03",X"1F",X"7C",
		X"E0",X"83",X"1F",X"78",X"F0",X"03",X"1F",X"7C",X"E0",X"83",X"1F",X"7C",X"F0",X"81",X"0F",X"7E",
		X"F0",X"C3",X"0F",X"7E",X"F0",X"83",X"1F",X"3E",X"F0",X"83",X"0F",X"7E",X"F0",X"83",X"1F",X"3E",
		X"F0",X"C3",X"07",X"7E",X"F8",X"C1",X"0F",X"7E",X"F0",X"C3",X"0B",X"7E",X"F8",X"C0",X"0F",X"3E",
		X"F0",X"C1",X"0F",X"7E",X"78",X"C1",X"0F",X"3E",X"F0",X"C3",X"03",X"7E",X"F0",X"81",X"1F",X"3E",
		X"E0",X"83",X"1F",X"7C",X"F0",X"03",X"1F",X"7C",X"E0",X"83",X"1F",X"F8",X"E0",X"07",X"3E",X"F8",
		X"C0",X"07",X"1F",X"F8",X"E0",X"07",X"3F",X"BC",X"E0",X"07",X"3F",X"F8",X"C1",X"07",X"3E",X"F8",
		X"C1",X"0F",X"1F",X"F8",X"C1",X"07",X"7E",X"78",X"C1",X"0F",X"3E",X"F8",X"C1",X"07",X"7E",X"F8",
		X"C0",X"0F",X"3E",X"F0",X"C3",X"0B",X"7E",X"F0",X"82",X"1F",X"3E",X"F0",X"83",X"0F",X"FC",X"F0",
		X"82",X"1F",X"FC",X"E0",X"87",X"17",X"FC",X"E0",X"07",X"3F",X"F8",X"C0",X"07",X"3F",X"F8",X"C1",
		X"07",X"7E",X"F0",X"81",X"1F",X"7E",X"E0",X"83",X"1F",X"F8",X"E0",X"07",X"3E",X"7C",X"C0",X"0F",
		X"2F",X"F0",X"C3",X"0B",X"FC",X"F0",X"01",X"3F",X"BC",X"C0",X"0F",X"1F",X"F0",X"83",X"0F",X"F8",
		X"E0",X"07",X"3E",X"7C",X"C0",X"0F",X"7E",X"E0",X"83",X"1F",X"F8",X"E0",X"07",X"3E",X"F8",X"01",
		X"1F",X"7E",X"C0",X"07",X"3F",X"F0",X"C1",X"1B",X"FC",X"E0",X"07",X"3E",X"DC",X"81",X"1F",X"D6",
		X"E0",X"07",X"3F",X"F0",X"C3",X"1B",X"F8",X"E0",X"07",X"7E",X"F0",X"03",X"3F",X"F8",X"81",X"1F",
		X"BC",X"C0",X"0F",X"7E",X"E0",X"83",X"37",X"F0",X"C1",X"17",X"F8",X"C1",X"1B",X"DC",X"E0",X"0F",
		X"FC",X"E0",X"06",X"7E",X"E0",X"07",X"7E",X"F0",X"06",X"6E",X"F0",X"06",X"7E",X"B0",X"07",X"7E",
		X"E0",X"07",X"5E",X"F0",X"03",X"DE",X"E0",X"05",X"BC",X"E0",X"1D",X"D8",X"C1",X"E9",X"30",X"C3",
		X"55",X"61",X"0E",X"1B",X"83",X"3D",X"0E",X"07",X"F3",X"B0",X"70",X"88",X"E3",X"A1",X"01",X"1F",
		X"8E",X"39",X"F0",X"F0",X"0C",X"1E",X"8A",X"07",X"FE",X"C0",X"F0",X"09",X"1E",X"16",X"CE",X"C2",
		X"07",X"CC",X"2F",X"E0",X"0B",X"F0",X"29",X"3E",X"70",X"F8",X"08",X"7E",X"02",X"F8",X"0F",X"26",
		X"71",X"2C",X"87",X"07",X"09",X"FF",X"80",X"3F",X"10",X"FE",X"03",X"EA",X"05",X"87",X"F0",X"03",
		X"1C",X"7F",X"00",X"7F",X"05",X"F8",X"07",X"62",X"3F",X"30",X"8E",X"0F",X"E0",X"7E",X"00",X"F7",
		X"71",X"E0",X"0F",X"1C",X"78",X"2E",X"02",X"3F",X"21",X"FC",X"09",X"E8",X"0F",X"38",X"87",X"0F",
		X"30",X"FE",X"00",X"7E",X"15",X"E5",X"38",X"CF",X"B1",X"AC",X"AA",X"AA",X"2A",X"55",X"55",X"55",
		X"10",X"CF",X"73",X"9C",X"AA",X"A6",X"CE",X"92",X"AD",X"8E",X"E5",X"54",X"65",X"CA",X"81",X"B1",
		X"98",X"D6",X"31",X"CB",X"D2",X"A6",X"2C",X"6B",X"59",X"5B",X"D2",X"B2",X"8C",X"66",X"6C",X"8C",
		X"18",X"E6",X"B4",X"8E",X"73",X"96",X"92",X"A7",X"9C",X"A6",X"32",X"C7",X"72",X"8E",X"69",X"CC",
		X"31",X"2B",X"33",X"B1",X"96",X"25",X"8D",X"69",X"0E",X"96",X"31",X"A5",X"31",X"9A",X"32",X"35",
		X"6C",X"98",X"51",X"32",X"53",X"72",X"39",X"76",X"7A",X"5A",X"5D",X"BC",X"3C",X"CE",X"39",X"CE",
		X"39",X"CF",X"BA",X"CE",X"AE",X"3D",X"D7",X"5E",X"37",X"C7",X"29",X"8E",X"E3",X"4C",X"87",X"73",
		X"C6",X"63",X"A5",X"CA",X"61",X"29",X"61",X"B1",X"54",X"65",X"34",X"A5",X"28",X"8C",X"54",X"51",
		X"51",X"A2",X"A2",X"35",X"D7",X"5C",X"AF",X"EB",X"6B",X"AF",X"B7",X"4D",X"AB",X"CE",X"B5",X"AD",
		X"AB",X"A6",X"21",X"C5",X"A4",X"88",X"29",X"12",X"21",X"09",X"92",X"90",X"A2",X"94",X"A2",X"44",
		X"45",X"B1",X"A2",X"95",X"5A",X"E9",X"6A",X"AD",X"54",X"55",X"5D",X"DD",X"B6",X"5E",X"B7",X"DF",
		X"DE",X"BE",X"DD",X"6E",X"B7",X"DB",X"ED",X"AE",X"AD",X"AD",X"B6",X"DA",X"5A",X"5D",X"D7",X"2E",
		X"AD",X"AA",X"10",X"0A",X"89",X"24",X"A9",X"A4",X"0A",X"95",X"54",X"45",X"55",X"6A",X"95",X"14",
		X"A9",X"64",X"49",X"51",X"51",X"25",X"51",X"4A",X"56",X"55",X"AA",X"2A",X"2A",X"54",X"89",X"12",
		X"94",X"94",X"2A",X"2A",X"A9",X"4A",X"55",X"55",X"D1",X"D2",X"55",X"69",X"D5",X"EB",X"AA",X"EB",
		X"D5",X"B7",X"DB",X"AB",X"D5",X"AA",X"D5",X"55",X"AB",X"45",X"95",X"B5",X"F5",X"AA",X"97",X"5B",
		X"ED",X"AA",X"B5",X"F4",X"52",X"2B",X"75",X"A8",X"52",X"A5",X"EA",X"B4",X"4B",X"48",X"10",X"41",
		X"20",X"48",X"50",X"28",X"B2",X"A8",X"AA",X"DA",X"7A",X"DD",X"DD",X"DD",X"F7",X"BD",X"BB",X"7D",
		X"DB",X"ED",X"AE",X"DA",X"6A",X"9B",X"A0",X"00",X"10",X"48",X"42",X"09",X"2A",X"50",X"49",X"5A",
		X"55",X"AB",X"56",X"77",X"BB",X"F7",X"7D",X"F7",X"BE",X"B7",X"B7",X"F7",X"DE",X"0E",X"05",X"14",
		X"44",X"14",X"24",X"44",X"88",X"24",X"A9",X"14",X"25",X"4A",X"95",X"AA",X"9A",X"57",X"AF",X"BB",
		X"D7",X"AF",X"DF",X"FD",X"76",X"B7",X"BB",X"D7",X"57",X"51",X"00",X"01",X"12",X"A1",X"04",X"09",
		X"92",X"88",X"2A",X"8A",X"8A",X"54",X"A5",X"56",X"B5",X"7A",X"DB",X"DD",X"FE",X"EE",X"77",X"EF",
		X"BE",X"FB",X"F6",X"DB",X"0E",X"03",X"02",X"85",X"0A",X"45",X"42",X"12",X"16",X"29",X"A5",X"94",
		X"A4",X"52",X"55",X"5A",X"B5",X"DB",X"ED",X"DD",X"7B",X"DF",X"BB",X"D7",X"DE",X"6E",X"6F",X"2B",
		X"0A",X"00",X"10",X"95",X"54",X"44",X"21",X"2A",X"A9",X"52",X"2A",X"52",X"A9",X"AA",X"5A",X"D5",
		X"57",X"AF",X"BE",X"76",X"BF",X"7B",X"7B",X"BB",X"BD",X"FA",X"5A",X"A1",X"00",X"80",X"40",X"91",
		X"22",X"42",X"42",X"91",X"AA",X"A4",X"92",X"AA",X"AA",X"75",X"B7",X"DB",X"ED",X"FB",X"F6",X"DB",
		X"EF",X"EF",X"DD",X"DE",X"EE",X"DA",X"AD",X"52",X"40",X"80",X"20",X"90",X"A0",X"90",X"48",X"A4",
		X"50",X"51",X"49",X"A5",X"52",X"A9",X"D5",X"5A",X"BB",X"F5",X"DA",X"DD",X"7E",X"EF",X"ED",X"EE",
		X"DD",X"56",X"57",X"AD",X"82",X"00",X"01",X"81",X"40",X"42",X"24",X"22",X"89",X"14",X"95",X"94",
		X"4A",X"55",X"AD",X"F5",X"DA",X"DB",X"BD",X"DE",X"BD",X"F7",X"B7",X"BB",X"FB",X"DA",X"6D",X"75",
		X"55",X"29",X"90",X"40",X"82",X"40",X"82",X"84",X"84",X"92",X"12",X"25",X"49",X"49",X"29",X"A5",
		X"54",X"55",X"ED",X"B6",X"BB",X"EF",X"7F",X"7F",X"BF",X"FB",X"FB",X"6E",X"AF",X"5E",X"55",X"05",
		X"25",X"28",X"20",X"02",X"04",X"22",X"88",X"08",X"09",X"49",X"A4",X"54",X"55",X"59",X"D5",X"DB",
		X"DD",X"FB",X"7E",X"FF",X"FD",X"EE",X"BB",X"EF",X"B6",X"6A",X"AA",X"14",X"44",X"00",X"01",X"81",
		X"08",X"12",X"22",X"91",X"24",X"A5",X"94",X"AA",X"AA",X"5A",X"AF",X"7B",X"FB",X"F6",X"DB",X"EF",
		X"FB",X"7B",X"D7",X"56",X"6B",X"B5",X"AA",X"24",X"11",X"20",X"40",X"20",X"88",X"20",X"44",X"22",
		X"51",X"54",X"A9",X"54",X"55",X"EB",X"D6",X"ED",X"ED",X"F6",X"FB",X"EB",X"75",X"75",X"F5",X"D6",
		X"6A",X"75",X"AD",X"55",X"55",X"1A",X"11",X"04",X"10",X"08",X"22",X"44",X"14",X"A5",X"94",X"4A",
		X"55",X"55",X"55",X"B7",X"5D",X"EF",X"D6",X"B6",X"5A",X"6D",X"75",X"EF",X"5D",X"BD",X"DE",X"6E",
		X"5B",X"97",X"8E",X"02",X"41",X"08",X"89",X"90",X"40",X"11",X"A5",X"54",X"A5",X"AA",X"AA",X"6A",
		X"EB",X"AA",X"45",X"D1",X"64",X"55",X"75",X"6D",X"7B",X"D7",X"BD",X"7B",X"5F",X"7B",X"5D",X"2B",
		X"12",X"A4",X"A0",X"90",X"44",X"92",X"A8",X"52",X"55",X"55",X"6A",X"55",X"75",X"D5",X"92",X"0A",
		X"16",X"8D",X"2A",X"AD",X"5E",X"BF",X"BE",X"DE",X"ED",X"F5",X"DA",X"AD",X"14",X"48",X"08",X"12",
		X"24",X"92",X"44",X"8A",X"2A",X"55",X"A9",X"AA",X"AA",X"AA",X"AA",X"53",X"15",X"2D",X"55",X"55",
		X"D5",X"7E",X"BD",X"BE",X"BE",X"DE",X"7A",X"AF",X"4A",X"10",X"44",X"02",X"85",X"22",X"45",X"8A",
		X"2A",X"55",X"55",X"D3",X"EA",X"D6",X"6D",X"5B",X"B7",X"5B",X"6B",X"ED",X"DA",X"76",X"BD",X"76",
		X"5D",X"5D",X"AF",X"AE",X"04",X"02",X"10",X"00",X"11",X"84",X"84",X"12",X"95",X"AA",X"AA",X"5A",
		X"D7",X"6E",X"6F",X"EF",X"DD",X"B7",X"77",X"BB",X"6D",X"5B",X"B7",X"5A",X"55",X"1A",X"34",X"A9",
		X"10",X"10",X"80",X"00",X"41",X"10",X"21",X"89",X"52",X"95",X"AA",X"56",X"BB",X"DE",X"EE",X"DE",
		X"BB",X"BF",X"77",X"BD",X"76",X"BD",X"B6",X"5A",X"B5",X"AA",X"AA",X"8A",X"0A",X"02",X"04",X"04",
		X"12",X"04",X"09",X"89",X"48",X"A5",X"2A",X"B5",X"AA",X"D6",X"75",X"D7",X"B7",X"AF",X"B7",X"DB",
		X"DB",X"DD",X"ED",X"DB",X"D5",X"56",X"D5",X"D2",X"42",X"85",X"80",X"00",X"80",X"10",X"42",X"44",
		X"44",X"92",X"54",X"AA",X"AA",X"AA",X"B6",X"DD",X"6D",X"B7",X"D7",X"F7",X"ED",X"DD",X"F7",X"BB",
		X"EF",X"AD",X"B7",X"B6",X"5A",X"B5",X"24",X"02",X"01",X"10",X"10",X"41",X"84",X"08",X"89",X"24",
		X"95",X"2A",X"55",X"AA",X"AA",X"AD",X"5D",X"6F",X"77",X"EF",X"BB",X"EF",X"EF",X"B7",X"AF",X"6F",
		X"77",X"B5",X"56",X"25",X"02",X"01",X"01",X"01",X"11",X"82",X"88",X"48",X"92",X"A4",X"A2",X"4A",
		X"55",X"55",X"55",X"AB",X"5B",X"6F",X"77",X"FB",X"FD",X"BE",X"EF",X"7D",X"F7",X"EE",X"AE",X"AD",
		X"2A",X"11",X"21",X"08",X"04",X"42",X"20",X"22",X"12",X"49",X"52",X"52",X"29",X"55",X"55",X"D5",
		X"EA",X"B6",X"ED",X"F6",X"EE",X"FB",X"F7",X"77",X"EF",X"B7",X"77",X"DB",X"D6",X"2A",X"25",X"10",
		X"10",X"40",X"10",X"04",X"21",X"44",X"24",X"49",X"4A",X"A5",X"2A",X"55",X"AD",X"6B",X"EB",X"B6",
		X"B7",X"DB",X"FB",X"FD",X"BB",X"6F",X"BF",X"DE",X"AE",X"AD",X"A6",X"82",X"10",X"02",X"02",X"81",
		X"20",X"42",X"44",X"24",X"49",X"52",X"A9",X"54",X"D5",X"6A",X"DD",X"76",X"7B",X"BB",X"DB",X"F7",
		X"FE",X"DE",X"DD",X"6F",X"6F",X"AF",X"AD",X"2A",X"05",X"08",X"10",X"20",X"40",X"08",X"21",X"24",
		X"51",X"51",X"29",X"55",X"D9",X"6A",X"DB",X"76",X"7B",X"F7",X"EE",X"EE",X"7D",X"DF",X"ED",X"F5",
		X"6D",X"DB",X"B6",X"55",X"05",X"02",X"01",X"40",X"80",X"80",X"10",X"44",X"22",X"49",X"52",X"AA",
		X"54",X"B5",X"DA",X"B6",X"BB",X"7D",X"DF",X"BE",X"6F",X"BF",X"DF",X"DD",X"BB",X"B7",X"DB",X"DA",
		X"AA",X"14",X"10",X"20",X"40",X"10",X"10",X"90",X"88",X"24",X"94",X"A4",X"92",X"AA",X"6A",X"D5",
		X"B5",X"BB",X"7D",X"F7",X"ED",X"F7",X"FE",X"BE",X"ED",X"ED",X"ED",X"DA",X"6A",X"91",X"80",X"00",
		X"01",X"01",X"10",X"84",X"10",X"91",X"48",X"A4",X"A4",X"52",X"55",X"55",X"B5",X"DB",X"BE",X"7D",
		X"F7",X"FE",X"FE",X"FE",X"EE",X"7E",X"F7",X"D6",X"AE",X"56",X"09",X"08",X"11",X"20",X"00",X"08",
		X"88",X"90",X"88",X"48",X"52",X"52",X"A9",X"54",X"B5",X"EA",X"76",X"FB",X"7B",X"DF",X"F7",X"BF",
		X"DF",X"7E",X"DF",X"DE",X"B6",X"AD",X"26",X"10",X"41",X"00",X"08",X"20",X"08",X"42",X"44",X"22",
		X"91",X"24",X"A9",X"4A",X"55",X"B5",X"AD",X"BB",X"7B",X"EF",X"FE",X"FD",X"FB",X"7B",X"BF",X"FB",
		X"AE",X"BD",X"25",X"11",X"22",X"02",X"00",X"01",X"21",X"84",X"88",X"24",X"89",X"24",X"A5",X"52",
		X"AA",X"6A",X"DD",X"B6",X"7D",X"DF",X"FB",X"FD",X"FD",X"7B",X"F7",X"77",X"6F",X"DB",X"2D",X"01",
		X"89",X"40",X"00",X"40",X"10",X"44",X"88",X"48",X"24",X"49",X"4A",X"AA",X"AA",X"D6",X"D6",X"6D",
		X"BF",X"DD",X"FB",X"FE",X"FB",X"BB",X"FD",X"77",X"6F",X"DB",X"2D",X"81",X"84",X"10",X"00",X"20",
		X"08",X"21",X"88",X"24",X"24",X"49",X"AA",X"A4",X"AA",X"DA",X"D6",X"76",X"FB",X"6E",X"EF",X"DF",
		X"EF",X"F7",X"7D",X"BF",X"DE",X"5B",X"BB",X"02",X"14",X"41",X"00",X"40",X"04",X"42",X"08",X"25",
		X"22",X"49",X"A9",X"52",X"5A",X"D5",X"B6",X"DD",X"DD",X"BD",X"FB",X"7B",X"FF",X"DD",X"FD",X"BD",
		X"7B",X"5B",X"B7",X"80",X"24",X"80",X"10",X"00",X"04",X"24",X"01",X"29",X"21",X"25",X"49",X"4B",
		X"55",X"55",X"7B",X"ED",X"DE",X"F6",X"B7",X"7F",X"F7",X"EF",X"DE",X"FD",X"EE",X"B6",X"5A",X"15",
		X"90",X"10",X"10",X"00",X"10",X"04",X"41",X"14",X"92",X"24",X"A5",X"54",X"55",X"D5",X"B6",X"DD",
		X"DD",X"7E",X"DF",X"77",X"7F",X"DF",X"BB",X"FB",X"5B",X"BB",X"AA",X"AA",X"00",X"21",X"10",X"00",
		X"10",X"84",X"40",X"14",X"91",X"24",X"A9",X"4A",X"AA",X"6A",X"BB",X"D6",X"7B",X"F7",X"FB",X"7E",
		X"DF",X"FB",X"DE",X"BD",X"BB",X"6D",X"55",X"55",X"0A",X"00",X"24",X"00",X"01",X"20",X"21",X"50",
		X"22",X"52",X"92",X"54",X"95",X"5A",X"F5",X"76",X"DD",X"FB",X"BE",X"F7",X"FE",X"DE",X"F7",X"EE",
		X"76",X"5B",X"55",X"55",X"89",X"20",X"00",X"21",X"00",X"80",X"10",X"21",X"24",X"A2",X"94",X"A4",
		X"AA",X"AC",X"AA",X"DE",X"6E",X"DF",X"FD",X"7B",X"EF",X"F7",X"BD",X"EF",X"AD",X"DD",X"AA",X"AA",
		X"92",X"14",X"04",X"10",X"02",X"02",X"10",X"12",X"42",X"92",X"50",X"4A",X"AA",X"4A",X"B5",X"5A",
		X"6F",X"FB",X"BE",X"F7",X"F7",X"BE",X"F7",X"BD",X"BB",X"D5",X"B6",X"4A",X"29",X"49",X"08",X"01",
		X"10",X"01",X"42",X"40",X"24",X"48",X"22",X"A5",X"94",X"AA",X"5A",X"55",X"6F",X"D7",X"F7",X"7B",
		X"7F",X"EF",X"77",X"F7",X"BB",X"55",X"6D",X"AB",X"52",X"45",X"89",X"20",X"10",X"10",X"20",X"10",
		X"08",X"49",X"44",X"4A",X"4A",X"95",X"AA",X"AA",X"75",X"DB",X"EE",X"F7",X"7D",X"EF",X"F7",X"BD",
		X"FB",X"5E",X"B5",X"D6",X"AA",X"52",X"52",X"12",X"08",X"40",X"02",X"10",X"04",X"A2",X"04",X"91",
		X"92",X"AA",X"52",X"B5",X"55",X"DD",X"DD",X"BD",X"7B",X"7F",X"EF",X"7B",X"F7",X"DE",X"AD",X"5A",
		X"AB",X"AA",X"12",X"A9",X"10",X"10",X"80",X"20",X"40",X"10",X"A2",X"10",X"29",X"A9",X"2A",X"55",
		X"AD",X"DA",X"B6",X"6F",X"EF",X"FB",X"7D",X"BF",X"F7",X"DE",X"BD",X"5B",X"ED",X"AA",X"5A",X"92",
		X"0A",X"10",X"80",X"08",X"00",X"82",X"10",X"11",X"49",X"92",X"52",X"95",X"5A",X"B5",X"AE",X"BD",
		X"BB",X"F7",X"FD",X"BB",X"F7",X"F7",X"EE",X"ED",X"EE",X"36",X"B5",X"55",X"A5",X"00",X"20",X"04",
		X"02",X"00",X"21",X"22",X"22",X"89",X"24",X"55",X"55",X"55",X"B5",X"76",X"77",X"77",X"EF",X"EF",
		X"7B",X"EF",X"EF",X"DD",X"DE",X"DE",X"55",X"B5",X"AA",X"12",X"00",X"12",X"00",X"02",X"40",X"12",
		X"90",X"24",X"52",X"92",X"AA",X"4A",X"AD",X"B6",X"BB",X"7D",X"FB",X"F7",X"DD",X"EF",X"FD",X"DE",
		X"BB",X"DD",X"DB",X"DA",X"AA",X"AA",X"04",X"40",X"00",X"01",X"00",X"11",X"84",X"48",X"44",X"91",
		X"54",X"AA",X"54",X"B5",X"6D",X"BB",X"FB",X"DE",X"F7",X"DD",X"BF",X"EF",X"BE",X"BB",X"77",X"B5",
		X"5B",X"55",X"05",X"88",X"04",X"08",X"00",X"48",X"80",X"48",X"88",X"14",X"51",X"AA",X"54",X"55",
		X"B5",X"DB",X"EE",X"DE",X"FB",X"DD",X"F7",X"FB",X"BE",X"EB",X"77",X"DB",X"B6",X"DA",X"92",X"40",
		X"04",X"08",X"00",X"10",X"02",X"89",X"10",X"89",X"A4",X"24",X"A9",X"52",X"B5",X"DA",X"DD",X"ED",
		X"FB",X"7D",X"EF",X"FD",X"7D",X"6F",X"F7",X"DB",X"76",X"AB",X"55",X"05",X"91",X"20",X"00",X"40",
		X"10",X"84",X"08",X"92",X"48",X"52",X"92",X"AA",X"54",X"6B",X"DD",X"6D",X"BF",X"FB",X"DD",X"F7",
		X"FB",X"BD",X"ED",X"77",X"B7",X"D5",X"5A",X"55",X"01",X"09",X"01",X"04",X"80",X"10",X"04",X"44",
		X"24",X"89",X"24",X"A5",X"AA",X"AA",X"B6",X"DB",X"EE",X"BD",X"DF",X"FD",X"BE",X"EF",X"BB",X"7B",
		X"EF",X"76",X"AD",X"B6",X"8A",X"40",X"21",X"10",X"00",X"42",X"10",X"11",X"24",X"22",X"29",X"49",
		X"95",X"AA",X"6A",X"DD",X"75",X"F7",X"EE",X"7D",X"F7",X"7B",X"7F",X"DB",X"7D",X"BB",X"5D",X"D5",
		X"2A",X"09",X"42",X"00",X"08",X"00",X"04",X"21",X"22",X"22",X"49",X"52",X"4A",X"55",X"55",X"EB",
		X"B6",X"77",X"EF",X"FD",X"BE",X"EF",X"7B",X"DF",X"DD",X"BB",X"DB",X"D6",X"56",X"15",X"21",X"04",
		X"04",X"40",X"00",X"11",X"44",X"44",X"24",X"91",X"92",X"AA",X"52",X"B5",X"DA",X"ED",X"EE",X"DE",
		X"FB",X"BE",X"EF",X"7D",X"6F",X"77",X"77",X"5B",X"AB",X"2A",X"45",X"10",X"08",X"10",X"10",X"10",
		X"22",X"24",X"12",X"25",X"49",X"95",X"AA",X"AA",X"5A",X"B7",X"DD",X"DD",X"7B",X"EF",X"DD",X"77",
		X"F7",X"EE",X"EE",X"DA",X"B6",X"55",X"55",X"89",X"04",X"41",X"08",X"20",X"04",X"21",X"22",X"92",
		X"48",X"4A",X"49",X"95",X"AA",X"AA",X"D6",X"6D",X"7B",X"EF",X"EE",X"DE",X"DE",X"DD",X"EE",X"6E",
		X"DB",X"56",X"55",X"15",X"09",X"04",X"11",X"40",X"10",X"44",X"44",X"24",X"29",X"49",X"29",X"55",
		X"55",X"55",X"AB",X"B7",X"DD",X"BD",X"F7",X"DD",X"BD",X"EF",X"F6",X"6E",X"77",X"6B",X"55",X"55",
		X"25",X"04",X"11",X"04",X"02",X"21",X"42",X"44",X"22",X"29",X"29",X"A9",X"54",X"55",X"D5",X"BA",
		X"DB",X"DD",X"7D",X"EF",X"DD",X"DD",X"BB",X"DB",X"DD",X"6E",X"5B",X"55",X"55",X"21",X"08",X"04",
		X"01",X"82",X"20",X"42",X"44",X"22",X"49",X"52",X"4A",X"A9",X"AA",X"6A",X"D7",X"ED",X"EE",X"BD",
		X"F7",X"EE",X"BE",X"7B",X"77",X"BB",X"DB",X"B6",X"AA",X"AA",X"84",X"10",X"08",X"01",X"81",X"20",
		X"42",X"44",X"22",X"49",X"4A",X"29",X"55",X"55",X"AD",X"DB",X"6D",X"EF",X"5D",X"DF",X"F7",X"EE",
		X"F7",X"DE",X"5D",X"B7",X"6D",X"55",X"55",X"22",X"21",X"10",X"80",X"20",X"10",X"22",X"44",X"12",
		X"49",X"49",X"A5",X"AA",X"AA",X"DA",X"DD",X"ED",X"BD",X"FB",X"DE",X"F7",X"DD",X"7D",X"77",X"B7",
		X"6E",X"AD",X"29",X"11",X"44",X"00",X"04",X"10",X"08",X"11",X"11",X"49",X"92",X"94",X"52",X"A5",
		X"AA",X"B5",X"DB",X"BB",X"EF",X"FD",X"BE",X"EF",X"7B",X"DF",X"7D",X"7B",X"BD",X"B5",X"AA",X"24",
		X"12",X"08",X"40",X"80",X"10",X"44",X"88",X"88",X"24",X"92",X"94",X"4A",X"55",X"D5",X"D6",X"DB",
		X"DE",X"BD",X"F7",X"FB",X"7D",X"BF",X"FB",X"EE",X"6E",X"5B",X"9A",X"12",X"11",X"01",X"04",X"82",
		X"20",X"82",X"88",X"88",X"48",X"92",X"54",X"4A",X"55",X"AD",X"76",X"BB",X"BB",X"7B",X"EF",X"EF",
		X"F7",X"7E",X"DF",X"BE",X"DB",X"96",X"26",X"15",X"21",X"02",X"44",X"88",X"10",X"11",X"12",X"22",
		X"22",X"12",X"25",X"A5",X"AA",X"AA",X"5A",X"B7",X"6D",X"77",X"FB",X"7E",X"DF",X"DF",X"DF",X"DE",
		X"DD",X"AA",X"AA",X"42",X"09",X"22",X"22",X"21",X"41",X"A2",X"90",X"90",X"88",X"48",X"92",X"94",
		X"AA",X"AA",X"6A",X"DD",X"B6",X"DD",X"FB",X"BE",X"F7",X"F7",X"F7",X"76",X"D7",X"53",X"93",X"8A",
		X"44",X"04",X"89",X"84",X"44",X"84",X"88",X"22",X"92",X"48",X"52",X"52",X"AA",X"AA",X"5A",X"B7",
		X"DB",X"DD",X"FB",X"DE",X"FB",X"D7",X"EF",X"EB",X"B5",X"55",X"A5",X"22",X"21",X"21",X"42",X"22",
		X"11",X"21",X"41",X"41",X"42",X"24",X"4A",X"52",X"4A",X"55",X"55",X"5B",X"B7",X"6E",X"DF",X"7B",
		X"F7",X"F7",X"F7",X"F6",X"BA",X"55",X"55",X"A9",X"28",X"21",X"11",X"89",X"48",X"24",X"11",X"11",
		X"91",X"44",X"12",X"29",X"A9",X"54",X"55",X"B5",X"7A",X"BB",X"F7",X"DE",X"FD",X"F6",X"DB",X"DD",
		X"76",X"DB",X"AA",X"24",X"49",X"22",X"41",X"22",X"22",X"21",X"91",X"48",X"88",X"48",X"48",X"12",
		X"29",X"A9",X"54",X"B5",X"D6",X"ED",X"EE",X"BD",X"F7",X"DD",X"DF",X"7E",X"7D",X"BB",X"6D",X"AD",
		X"AA",X"54",X"41",X"85",X"44",X"22",X"84",X"04",X"11",X"08",X"21",X"22",X"91",X"A2",X"54",X"55",
		X"D5",X"D6",X"DB",X"DD",X"FD",X"BE",X"F7",X"FD",X"BE",X"77",X"B7",X"5D",X"6B",X"55",X"A5",X"8A",
		X"24",X"11",X"41",X"02",X"81",X"10",X"08",X"04",X"09",X"49",X"94",X"4A",X"55",X"55",X"BB",X"6E",
		X"77",X"77",X"EF",X"7D",X"DF",X"BB",X"B7",X"77",X"D7",X"56",X"55",X"2A",X"49",X"12",X"22",X"04",
		X"11",X"10",X"04",X"02",X"11",X"92",X"88",X"2A",X"55",X"D5",X"DA",X"ED",X"DE",X"7D",X"BF",X"EF",
		X"BD",X"DF",X"77",X"F7",X"76",X"5B",X"55",X"55",X"2A",X"52",X"88",X"90",X"10",X"04",X"11",X"88",
		X"10",X"22",X"89",X"24",X"95",X"AA",X"5A",X"AD",X"DD",X"DE",X"7B",X"BF",X"FB",X"FB",X"EE",X"BD",
		X"BB",X"5D",X"D5",X"4A",X"45",X"49",X"24",X"84",X"20",X"44",X"08",X"11",X"24",X"24",X"12",X"29",
		X"A5",X"52",X"55",X"6D",X"BD",X"EE",X"DE",X"F7",X"BE",X"DF",X"7B",X"EF",X"EE",X"ED",X"AA",X"95",
		X"2A",X"52",X"24",X"21",X"42",X"44",X"04",X"21",X"42",X"44",X"44",X"A2",X"92",X"4A",X"55",X"B5",
		X"76",X"DB",X"DD",X"F7",X"7D",X"DF",X"F7",X"7B",X"EF",X"DD",X"6D",X"5A",X"AA",X"28",X"22",X"11",
		X"11",X"12",X"12",X"11",X"22",X"22",X"12",X"91",X"24",X"A5",X"52",X"55",X"B5",X"DE",X"76",X"7B",
		X"DF",X"EF",X"DF",X"F7",X"7D",X"F7",X"DD",X"AA",X"52",X"45",X"12",X"11",X"89",X"48",X"48",X"50",
		X"44",X"42",X"88",X"88",X"24",X"25",X"95",X"AA",X"6A",X"B5",X"DB",X"75",X"EF",X"77",X"DF",X"F7",
		X"FB",X"BE",X"BD",X"55",X"95",X"92",X"44",X"42",X"42",X"12",X"49",X"24",X"91",X"88",X"48",X"24",
		X"92",X"92",X"4A",X"55",X"D5",X"D5",X"EB",X"D5",X"EB",X"BB",X"6F",X"BF",X"BF",X"7E",X"B7",X"AD",
		X"2A",X"29",X"14",X"51",X"28",X"49",X"52",X"4A",X"92",X"48",X"21",X"11",X"91",X"24",X"49",X"45",
		X"95",X"AA",X"AA",X"D5",X"ED",X"7D",X"F7",X"FE",X"FD",X"EE",X"DD",X"AB",X"AA",X"54",X"24",X"85",
		X"8A",X"2A",X"AA",X"54",X"4A",X"25",X"11",X"89",X"48",X"A2",X"28",X"49",X"A9",X"A8",X"2A",X"55",
		X"D5",X"D6",X"6F",X"BF",X"FD",X"7D",X"7B",X"BB",X"5A",X"A5",X"22",X"89",X"12",X"45",X"49",X"45",
		X"55",X"A5",X"A4",X"90",X"42",X"25",X"49",X"92",X"54",X"52",X"A5",X"52",X"D5",X"B6",X"DF",X"DB",
		X"DF",X"F7",X"BE",X"BB",X"DB",X"6A",X"A9",X"52",X"49",X"49",X"A9",X"A4",X"52",X"A9",X"52",X"51",
		X"44",X"A4",X"90",X"24",X"91",X"54",X"52",X"AA",X"D4",X"D2",X"D5",X"F7",X"7A",X"DB",X"B7",X"6F",
		X"77",X"55",X"95",X"42",X"49",X"8A",X"92",X"52",X"A5",X"52",X"55",X"55",X"92",X"48",X"48",X"24",
		X"45",X"8A",X"4A",X"95",X"AA",X"AA",X"AE",X"77",X"BD",X"FD",X"BE",X"7D",X"DD",X"B6",X"AA",X"4A",
		X"51",X"49",X"A5",X"54",X"55",X"55",X"D5",X"6E",X"AD",X"12",X"49",X"94",X"94",X"4A",X"94",X"94",
		X"2A",X"95",X"5A",X"5D",X"5F",X"AF",X"6F",X"6F",X"6F",X"57",X"97",X"4A",X"24",X"22",X"49",X"51",
		X"D1",X"D2",X"AA",X"D5",X"D5",X"2A",X"95",X"54",X"54",X"A4",X"A4",X"54",X"52",X"4A",X"55",X"AA",
		X"BA",X"7A",X"77",X"BD",X"AE",X"9E",X"2A",X"44",X"42",X"82",X"22",X"29",X"55",X"B5",X"FA",X"76",
		X"BB",X"BD",X"6D",X"AD",X"B6",X"AA",X"AA",X"56",X"95",X"2A",X"AB",X"AE",X"AD",X"D6",X"D6",X"D5",
		X"AB",X"25",X"41",X"10",X"90",X"20",X"21",X"51",X"4A",X"55",X"B5",X"D6",X"DB",X"6D",X"B7",X"DB",
		X"AE",X"6D",X"DB",X"DA",X"DA",X"DA",X"6A",X"D5",X"56",X"AB",X"AB",X"AE",X"2A",X"41",X"20",X"01",
		X"81",X"90",X"50",X"52",X"A5",X"AA",X"5A",X"7B",X"DD",X"76",X"7B",X"BB",X"DD",X"7A",X"B5",X"D5",
		X"AA",X"AA",X"4A",X"54",X"49",X"4A",X"55",X"4A",X"25",X"0A",X"08",X"08",X"08",X"11",X"45",X"A5",
		X"AA",X"AA",X"5A",X"77",X"DB",X"ED",X"EE",X"ED",X"ED",X"DB",X"B5",X"6D",X"AD",X"AA",X"AA",X"A8",
		X"28",X"A5",X"94",X"94",X"24",X"89",X"44",X"44",X"24",X"92",X"24",X"55",X"55",X"55",X"6D",X"7D",
		X"7B",X"BB",X"77",X"77",X"77",X"BB",X"DD",X"B6",X"5A",X"55",X"15",X"25",X"49",X"52",X"22",X"49",
		X"92",X"22",X"89",X"12",X"25",X"49",X"92",X"44",X"A5",X"54",X"95",X"AA",X"B6",X"F6",X"ED",X"F6",
		X"76",X"B7",X"BB",X"DB",X"AE",X"D6",X"AA",X"2A",X"52",X"14",X"25",X"45",X"49",X"49",X"29",X"29",
		X"49",X"52",X"92",X"24",X"A5",X"AA",X"AA",X"6A",X"6B",X"EF",X"ED",X"EE",X"B6",X"B7",X"DB",X"EE",
		X"76",X"6B",X"AD",X"AA",X"8A",X"24",X"91",X"24",X"89",X"24",X"4A",X"29",X"49",X"49",X"4A",X"92",
		X"A4",X"92",X"4A",X"55",X"D5",X"EA",X"EA",X"DB",X"5D",X"B7",X"7B",X"DD",X"76",X"DB",X"B6",X"B5",
		X"AA",X"8A",X"12",X"25",X"92",X"92",X"24",X"25",X"95",X"4A",X"4A",X"92",X"92",X"A8",X"54",X"51",
		X"55",X"55",X"D5",X"AA",X"F5",X"DD",X"D6",X"EB",X"AD",X"DB",X"36",X"5E",X"57",X"55",X"45",X"45",
		X"89",X"92",X"A4",X"94",X"52",X"A5",X"4A",X"55",X"95",X"54",X"4A",X"45",X"55",X"55",X"D5",X"AA",
		X"AB",X"D3",X"5D",X"D7",X"D6",X"6B",X"5B",X"DB",X"55",X"55",X"52",X"28",X"14",X"25",X"8C",X"62",
		X"A9",X"D4",X"B8",X"AA",X"E6",X"72",X"39",X"AE",X"55",X"3C",X"4D",X"E5",X"1C",X"C7",X"79",X"1E",
		X"8F",X"F3",X"B8",X"9C",X"2E",X"8B",X"59",X"52",X"C5",X"68",X"14",X"95",X"4C",X"1C",X"8E",X"D3",
		X"54",X"1E",X"9B",X"69",X"96",X"9A",X"2E",X"C7",X"99",X"CD",X"31",X"E7",X"CC",X"E3",X"32",X"C7",
		X"E3",X"70",X"98",X"C3",X"70",X"8C",X"D1",X"68",X"64",X"71",X"9A",X"E6",X"62",X"1E",X"9E",X"C7",
		X"B3",X"5A",X"66",X"73",X"35",X"CB",X"9A",X"99",X"1C",X"3C",X"8E",X"63",X"8E",X"C6",X"91",X"C1",
		X"61",X"12",X"C7",X"C8",X"98",X"C9",X"69",X"9A",X"CB",X"63",X"33",X"CF",X"A9",X"E3",X"99",X"73",
		X"E5",X"E3",X"B1",X"6A",X"78",X"78",X"78",X"38",X"3A",X"B1",X"4C",X"5C",X"3A",X"1C",X"6D",X"2C",
		X"36",X"3C",X"4E",X"79",X"64",X"39",X"76",X"5C",X"B5",X"5C",X"1C",X"D7",X"D1",X"46",X"8B",X"95",
		X"5A",X"1C",X"56",X"39",X"AA",X"72",X"D4",X"E2",X"61",X"C5",X"C5",X"99",X"8D",X"25",X"1E",X"8E",
		X"35",X"1E",X"8F",X"2B",X"17",X"4F",X"75",X"3A",X"1D",X"97",X"2E",X"9A",X"A9",X"AA",X"32",X"A5",
		X"CA",X"92",X"16",X"53",X"A5",X"91",X"C3",X"38",X"49",X"33",X"1E",X"2D",X"8D",X"8F",X"8B",X"47",
		X"37",X"6B",X"95",X"87",X"C7",X"CA",X"C3",X"A3",X"51",X"55",X"71",X"4C",X"55",X"9A",X"AA",X"9A",
		X"4A",X"39",X"AE",X"6C",X"7C",X"3C",X"3D",X"79",X"3C",X"AE",X"3A",X"3C",X"3C",X"38",X"38",X"18",
		X"1A",X"3A",X"5C",X"5C",X"5A",X"2E",X"6D",X"3A",X"AA",X"EA",X"74",X"75",X"F3",X"79",X"F5",X"F4",
		X"5A",X"1A",X"28",X"50",X"20",X"51",X"34",X"B5",X"F2",X"68",X"55",X"55",X"5A",X"CA",X"A2",X"51",
		X"0E",X"57",X"BD",X"AE",X"B7",X"AF",X"B7",X"DD",X"6E",X"DF",X"AE",X"47",X"05",X"0A",X"04",X"12",
		X"95",X"4A",X"AB",X"AA",X"AA",X"52",X"4A",X"11",X"4A",X"54",X"6A",X"F9",X"F5",X"ED",X"ED",X"7A",
		X"DD",X"DE",X"7B",X"78",X"30",X"A0",X"80",X"08",X"55",X"6A",X"59",X"55",X"2D",X"35",X"AA",X"54",
		X"0A",X"87",X"16",X"8F",X"77",X"BD",X"DB",X"ED",X"F5",X"7A",X"BD",X"7D",X"1B",X"0F",X"05",X"04",
		X"90",X"90",X"4A",X"55",X"AD",X"AA",X"AA",X"52",X"A5",X"42",X"45",X"A9",X"54",X"DB",X"BB",X"7B",
		X"EF",X"5E",X"AF",X"EB",X"5E",X"EF",X"E9",X"42",X"01",X"01",X"42",X"88",X"D2",X"34",X"CB",X"65",
		X"55",X"55",X"49",X"52",X"4A",X"49",X"AD",X"76",X"F7",X"DD",X"AE",X"B7",X"6D",X"F7",X"EC",X"F5",
		X"E9",X"60",X"40",X"80",X"20",X"48",X"B4",X"54",X"55",X"B5",X"CA",X"52",X"A9",X"A4",X"52",X"AA",
		X"5C",X"BD",X"DB",X"D7",X"5B",X"D7",X"AB",X"EB",X"F5",X"FA",X"E5",X"C3",X"08",X"01",X"41",X"88",
		X"B0",X"54",X"AA",X"6A",X"6A",X"2C",X"55",X"32",X"15",X"53",X"D5",X"BA",X"BB",X"DD",X"5E",X"AF",
		X"CE",X"6B",X"D7",X"EE",X"BE",X"3C",X"2C",X"10",X"10",X"08",X"12",X"8E",X"2A",X"4B",X"AB",X"CA",
		X"52",X"A5",X"4A",X"69",X"E9",X"F4",X"76",X"B7",X"BB",X"6E",X"5D",X"3D",X"5B",X"AF",X"7D",X"7D",
		X"79",X"18",X"10",X"10",X"10",X"11",X"15",X"4B",X"95",X"96",X"AA",X"52",X"A5",X"52",X"A9",X"B2",
		X"7C",X"7A",X"5D",X"D7",X"B5",X"AE",X"B5",X"AE",X"DB",X"DD",X"5B",X"3D",X"0C",X"08",X"04",X"82",
		X"42",X"A5",X"54",X"65",X"A9",X"52",X"32",X"54",X"28",X"4A",X"AA",X"AA",X"ED",X"EB",X"6E",X"B7",
		X"75",X"D7",X"DD",X"77",X"BF",X"3F",X"1D",X"2B",X"08",X"04",X"20",X"84",X"A2",X"52",X"95",X"AA",
		X"52",X"A9",X"94",X"54",X"52",X"55",X"D5",X"DB",X"BB",X"7B",X"7B",X"BB",X"DB",X"DB",X"FB",X"FD",
		X"3D",X"1E",X"06",X"08",X"80",X"20",X"12",X"A5",X"52",X"95",X"2A",X"A5",X"A4",X"24",X"49",X"A5",
		X"AA",X"ED",X"7D",X"F7",X"DE",X"DD",X"5B",X"CF",X"2B",X"57",X"57",X"57",X"0E",X"0A",X"04",X"20",
		X"20",X"91",X"A2",X"52",X"55",X"A5",X"2A",X"4D",X"55",X"55",X"D5",X"B5",X"D7",X"F7",X"BD",X"5B",
		X"57",X"2D",X"55",X"29",X"A7",X"DE",X"5D",X"35",X"14",X"10",X"00",X"04",X"11",X"45",X"55",X"55",
		X"B3",X"AA",X"55",X"4D",X"B5",X"5A",X"BB",X"BD",X"F3",X"EA",X"AA",X"AA",X"AA",X"D4",X"E6",X"B5",
		X"77",X"DF",X"D5",X"50",X"80",X"00",X"10",X"12",X"A9",X"54",X"B5",X"56",X"55",X"55",X"D5",X"72",
		X"A9",X"E3",X"4A",X"55",X"55",X"D5",X"71",X"D5",X"D5",X"5D",X"77",X"7D",X"7D",X"AD",X"06",X"09",
		X"04",X"80",X"90",X"A4",X"54",X"55",X"55",X"B5",X"AA",X"2E",X"2D",X"AA",X"54",X"2A",X"55",X"56",
		X"B5",X"EB",X"CE",X"EB",X"EA",X"79",X"ED",X"ED",X"36",X"1D",X"24",X"08",X"08",X"42",X"A2",X"92",
		X"A5",X"96",X"55",X"AD",X"3A",X"AA",X"54",X"14",X"A5",X"8A",X"AB",X"5E",X"AF",X"EB",X"D6",X"75",
		X"EB",X"F5",X"7A",X"6F",X"6D",X"9A",X"20",X"08",X"22",X"12",X"A5",X"52",X"55",X"CB",X"69",X"8E",
		X"52",X"14",X"12",X"49",X"4A",X"55",X"AD",X"BB",X"6E",X"5B",X"DB",X"5A",X"AF",X"DD",X"DB",X"4E",
		X"A3",X"00",X"81",X"20",X"24",X"A9",X"54",X"59",X"D5",X"9A",X"A6",X"8A",X"92",X"28",X"54",X"54",
		X"B5",X"EE",X"5E",X"D7",X"AE",X"D5",X"D6",X"D6",X"AD",X"B7",X"D7",X"3A",X"2A",X"20",X"08",X"91",
		X"94",X"4A",X"AD",X"D5",X"6B",X"D3",X"92",X"44",X"88",X"84",X"12",X"95",X"D5",X"7A",X"D7",X"75",
		X"6D",X"6D",X"ED",X"7A",X"DD",X"B6",X"5D",X"8D",X"0A",X"04",X"11",X"91",X"52",X"55",X"6B",X"B7",
		X"16",X"23",X"22",X"84",X"50",X"A2",X"52",X"B5",X"F5",X"B6",X"5D",X"D7",X"56",X"D7",X"BA",X"ED",
		X"7D",X"BB",X"EB",X"AA",X"28",X"28",X"24",X"24",X"54",X"54",X"AA",X"D2",X"A8",X"44",X"21",X"21",
		X"24",X"49",X"95",X"56",X"EB",X"6E",X"D7",X"DB",X"6E",X"D7",X"F7",X"FA",X"FA",X"BA",X"5A",X"45",
		X"44",X"08",X"44",X"44",X"49",X"55",X"AA",X"AA",X"A9",X"92",X"22",X"51",X"28",X"A9",X"AA",X"ED",
		X"BB",X"BD",X"BB",X"DB",X"DD",X"76",X"DB",X"DD",X"ED",X"6A",X"29",X"10",X"08",X"42",X"48",X"94",
		X"4A",X"55",X"55",X"35",X"55",X"2A",X"14",X"89",X"22",X"A5",X"AA",X"B5",X"77",X"BB",X"DB",X"AD",
		X"D7",X"DB",X"ED",X"D6",X"D5",X"4A",X"21",X"84",X"20",X"84",X"44",X"4A",X"95",X"AA",X"D5",X"DA",
		X"D2",X"51",X"45",X"49",X"92",X"4A",X"55",X"5D",X"6F",X"AF",X"77",X"B7",X"B7",X"DB",X"75",X"6B",
		X"55",X"29",X"10",X"41",X"10",X"91",X"28",X"A9",X"54",X"55",X"D5",X"EA",X"B2",X"56",X"AA",X"34",
		X"55",X"55",X"AD",X"5E",X"BB",X"DB",X"76",X"DB",X"EB",X"D5",X"B5",X"D6",X"52",X"40",X"40",X"20",
		X"48",X"A4",X"94",X"AA",X"AA",X"AA",X"AA",X"6B",X"6D",X"6B",X"EB",X"6A",X"6B",X"6D",X"6D",X"DB",
		X"75",X"BD",X"B6",X"7B",X"BB",X"EB",X"56",X"95",X"02",X"01",X"80",X"40",X"08",X"25",X"55",X"AA",
		X"4A",X"55",X"55",X"55",X"AD",X"DA",X"BA",X"BA",X"B6",X"75",X"ED",X"DA",X"DA",X"BA",X"B6",X"BD",
		X"D7",X"5D",X"5B",X"25",X"10",X"00",X"20",X"10",X"A2",X"94",X"52",X"55",X"55",X"55",X"55",X"55",
		X"D5",X"B6",X"DD",X"BE",X"DE",X"6E",X"D7",X"D6",X"5A",X"6D",X"75",X"BD",X"DD",X"6E",X"D5",X"04",
		X"02",X"20",X"80",X"20",X"92",X"54",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"BA",X"B6",X"BB",
		X"B7",X"5D",X"BB",X"56",X"6B",X"AD",X"75",X"B7",X"AF",X"3B",X"2D",X"05",X"02",X"08",X"10",X"84",
		X"44",X"49",X"A5",X"AA",X"AA",X"6A",X"55",X"B5",X"B6",X"AE",X"BB",X"DD",X"BB",X"DD",X"B6",X"55",
		X"AD",X"AA",X"34",X"AA",X"5A",X"55",X"22",X"10",X"10",X"00",X"08",X"42",X"24",X"29",X"55",X"A5",
		X"56",X"B5",X"BA",X"B6",X"DD",X"DE",X"DD",X"77",X"EF",X"76",X"5B",X"AB",X"55",X"55",X"55",X"D5",
		X"6A",X"55",X"4A",X"08",X"04",X"04",X"02",X"21",X"A2",X"A4",X"54",X"55",X"D5",X"EA",X"5A",X"6B",
		X"DB",X"B6",X"B7",X"6F",X"B7",X"DB",X"DA",X"AA",X"AA",X"AA",X"54",X"55",X"DD",X"AA",X"50",X"10",
		X"10",X"08",X"10",X"84",X"44",X"29",X"95",X"AA",X"6A",X"B5",X"BA",X"B5",X"ED",X"76",X"B7",X"B7",
		X"D7",X"6D",X"6B",X"6B",X"55",X"B5",X"5A",X"B5",X"5A",X"55",X"42",X"02",X"02",X"22",X"08",X"91",
		X"50",X"52",X"A9",X"AA",X"AA",X"75",X"DB",X"6E",X"77",X"EF",X"EE",X"F6",X"BA",X"6D",X"5B",X"AD",
		X"96",X"AA",X"94",X"AA",X"4A",X"45",X"42",X"10",X"08",X"02",X"21",X"12",X"49",X"52",X"AA",X"AA",
		X"6A",X"D5",X"6B",X"DB",X"F6",X"F6",X"F6",X"76",X"BB",X"75",X"B5",X"AA",X"AA",X"5A",X"AD",X"B6",
		X"5A",X"55",X"50",X"24",X"08",X"21",X"22",X"44",X"92",X"94",X"AA",X"54",X"D5",X"5A",X"F5",X"76",
		X"BB",X"7B",X"BB",X"EB",X"D6",X"55",X"AB",X"AA",X"94",X"54",X"A9",X"54",X"55",X"14",X"12",X"82",
		X"04",X"41",X"22",X"A2",X"24",X"A9",X"54",X"55",X"B5",X"BA",X"6E",X"7D",X"BD",X"7D",X"77",X"BB",
		X"5D",X"6B",X"AB",X"55",X"55",X"AD",X"56",X"5B",X"5B",X"55",X"21",X"84",X"20",X"21",X"91",X"48",
		X"51",X"A9",X"54",X"55",X"AA",X"AA",X"56",X"ED",X"ED",X"ED",X"BD",X"DD",X"B6",X"5A",X"AD",X"2A",
		X"AA",X"4A",X"4D",X"47",X"8F",X"8B",X"12",X"11",X"21",X"84",X"10",X"91",X"A4",X"92",X"2A",X"55",
		X"55",X"55",X"AB",X"B7",X"DB",X"BB",X"EF",X"76",X"B7",X"AD",X"55",X"AB",X"55",X"B5",X"EA",X"EA",
		X"DA",X"6A",X"55",X"08",X"09",X"22",X"44",X"24",X"49",X"25",X"55",X"95",X"AA",X"AA",X"AA",X"AA",
		X"6A",X"EF",X"76",X"B7",X"6B",X"5B",X"B5",X"AA",X"4A",X"A9",X"AC",X"5A",X"5A",X"AA",X"24",X"01",
		X"82",X"20",X"21",X"51",X"51",X"55",X"B5",X"6A",X"75",X"A9",X"AA",X"AA",X"6B",X"DB",X"DB",X"DD",
		X"DB",X"B6",X"AD",X"56",X"95",X"54",X"55",X"59",X"55",X"55",X"49",X"84",X"80",X"10",X"21",X"12",
		X"29",X"A9",X"AA",X"6A",X"55",X"AB",X"AA",X"6B",X"B7",X"B7",X"EF",X"BD",X"DB",X"ED",X"DA",X"AA",
		X"55",X"A5",X"54",X"A9",X"54",X"29",X"49",X"10",X"08",X"21",X"84",X"24",X"49",X"45",X"55",X"55",
		X"AD",X"BA",X"D6",X"BA",X"7A",X"DD",X"DD",X"BD",X"BB",X"B7",X"DB",X"B6",X"D5",X"6A",X"55",X"AD",
		X"AA",X"14",X"45",X"44",X"08",X"12",X"42",X"22",X"49",X"49",X"95",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"6A",X"6F",X"77",X"AF",X"77",X"B7",X"6B",X"5B",X"B5",X"AA",X"AA",X"92",X"AA",X"14",X"89",X"40",
		X"84",X"04",X"09",X"49",X"52",X"AA",X"54",X"D5",X"6A",X"75",X"6D",X"6B",X"BB",X"DD",X"BD",X"7B",
		X"EF",X"EE",X"6E",X"BB",X"56",X"5B",X"6D",X"5A",X"55",X"24",X"11",X"84",X"10",X"84",X"90",X"48",
		X"92",X"52",X"55",X"55",X"D5",X"EA",X"D2",X"D5",X"DA",X"76",X"BB",X"77",X"EF",X"EE",X"76",X"BB",
		X"BA",X"DA",X"AA",X"AA",X"4A",X"91",X"10",X"41",X"04",X"21",X"42",X"44",X"92",X"94",X"54",X"AA",
		X"AA",X"AA",X"6A",X"75",X"6D",X"BB",X"ED",X"DE",X"7B",X"77",X"F7",X"B6",X"EB",X"DA",X"EA",X"AA",
		X"A5",X"45",X"0A",X"09",X"11",X"44",X"10",X"11",X"11",X"49",X"29",X"55",X"55",X"55",X"55",X"AD",
		X"BA",X"B6",X"DD",X"DD",X"BB",X"77",X"F7",X"76",X"DB",X"75",X"B5",X"6A",X"55",X"15",X"09",X"09",
		X"02",X"09",X"44",X"88",X"48",X"A2",X"A4",X"4A",X"55",X"55",X"AB",X"DA",X"D6",X"B6",X"DD",X"DE",
		X"DD",X"BB",X"7B",X"EF",X"DD",X"6D",X"B7",X"B6",X"5A",X"55",X"15",X"49",X"08",X"11",X"84",X"10",
		X"12",X"91",X"24",X"49",X"A9",X"54",X"55",X"95",X"AA",X"AA",X"56",X"6F",X"B7",X"7D",X"7B",X"77",
		X"B7",X"EB",X"D6",X"56",X"AB",X"AA",X"28",X"91",X"40",X"10",X"41",X"44",X"48",X"24",X"49",X"52",
		X"A9",X"AA",X"AA",X"6A",X"F5",X"BA",X"6D",X"BB",X"BB",X"77",X"77",X"F7",X"7A",X"DB",X"75",X"6D",
		X"D5",X"52",X"51",X"22",X"44",X"10",X"42",X"08",X"11",X"49",X"92",X"94",X"4A",X"55",X"55",X"AB",
		X"6B",X"EB",X"B6",X"BD",X"DD",X"DD",X"DD",X"EE",X"76",X"DB",X"5D",X"5B",X"AB",X"56",X"85",X"44",
		X"04",X"09",X"42",X"88",X"88",X"24",X"49",X"49",X"95",X"AA",X"AA",X"AA",X"75",X"DB",X"DE",X"76",
		X"77",X"7B",X"BB",X"DD",X"5E",X"B7",X"AE",X"D5",X"6A",X"55",X"45",X"11",X"41",X"08",X"21",X"44",
		X"44",X"44",X"92",X"94",X"54",X"AA",X"54",X"55",X"D5",X"B6",X"DB",X"ED",X"76",X"B7",X"B7",X"B7",
		X"BD",X"5E",X"DB",X"D6",X"56",X"AB",X"8A",X"42",X"42",X"10",X"84",X"20",X"42",X"22",X"49",X"52",
		X"2A",X"A9",X"AA",X"AA",X"6A",X"DD",X"6E",X"6F",X"6F",X"6F",X"77",X"7B",X"BB",X"6D",X"DB",X"56",
		X"57",X"AD",X"2A",X"12",X"41",X"08",X"82",X"08",X"11",X"49",X"52",X"52",X"52",X"55",X"55",X"55",
		X"BB",X"ED",X"76",X"77",X"EF",X"EE",X"6E",X"77",X"DB",X"B6",X"D5",X"D5",X"AA",X"4A",X"11",X"21",
		X"02",X"81",X"10",X"42",X"44",X"92",X"A4",X"A4",X"52",X"55",X"55",X"D5",X"EA",X"6D",X"77",X"77",
		X"77",X"77",X"7B",X"DD",X"B6",X"AD",X"55",X"57",X"55",X"15",X"89",X"10",X"82",X"20",X"84",X"48",
		X"22",X"49",X"A5",X"54",X"55",X"55",X"55",X"B5",X"6E",X"B7",X"BB",X"BB",X"DB",X"DD",X"B6",X"6D",
		X"DB",X"DA",X"5A",X"B5",X"AA",X"8A",X"92",X"88",X"10",X"11",X"12",X"91",X"48",X"92",X"A4",X"94",
		X"52",X"A5",X"AA",X"AA",X"6A",X"ED",X"ED",X"EE",X"F6",X"6E",X"B7",X"DB",X"B6",X"AD",X"B5",X"56",
		X"55",X"95",X"14",X"45",X"84",X"10",X"22",X"88",X"88",X"44",X"92",X"A4",X"A4",X"52",X"A5",X"AA",
		X"AA",X"6A",X"BD",X"DD",X"DD",X"ED",X"76",X"DB",X"6D",X"DB",X"B6",X"B6",X"B5",X"6A",X"55",X"91",
		X"84",X"08",X"41",X"44",X"24",X"92",X"A4",X"94",X"52",X"95",X"AA",X"AA",X"AA",X"5A",X"6F",X"77",
		X"F7",X"F6",X"F6",X"76",X"DB",X"B6",X"6D",X"6D",X"D5",X"AA",X"AA",X"50",X"22",X"44",X"10",X"11",
		X"22",X"22",X"49",X"52",X"4A",X"A5",X"AA",X"AA",X"AA",X"AA",X"D6",X"DB",X"6E",X"77",X"77",X"BB",
		X"DD",X"B6",X"6D",X"6D",X"B5",X"6A",X"55",X"45",X"12",X"11",X"22",X"88",X"88",X"48",X"A4",X"24",
		X"A9",X"54",X"AA",X"54",X"55",X"AD",X"D6",X"DB",X"DD",X"DD",X"DD",X"ED",X"76",X"DB",X"76",X"6B",
		X"DB",X"6A",X"AD",X"AA",X"48",X"44",X"08",X"21",X"42",X"08",X"89",X"24",X"29",X"49",X"A5",X"52",
		X"95",X"AA",X"AA",X"B6",X"DE",X"EE",X"76",X"77",X"BB",X"BB",X"DD",X"6E",X"B7",X"5B",X"D7",X"6A",
		X"95",X"42",X"44",X"10",X"11",X"91",X"44",X"49",X"49",X"A5",X"4A",X"A9",X"52",X"A9",X"AA",X"AA",
		X"DD",X"DD",X"6E",X"B7",X"DD",X"DD",X"6E",X"B7",X"DD",X"B6",X"AB",X"55",X"15",X"12",X"84",X"10",
		X"41",X"44",X"24",X"49",X"92",X"92",X"54",X"2A",X"55",X"A9",X"AA",X"7A",X"7B",X"77",X"EF",X"EE",
		X"EE",X"5E",X"6F",X"BB",X"5D",X"B7",X"B6",X"2A",X"21",X"08",X"01",X"02",X"84",X"10",X"89",X"94",
		X"24",X"A5",X"52",X"A9",X"AA",X"6A",X"DD",X"ED",X"BB",X"EF",X"DB",X"77",X"F7",X"EE",X"ED",X"EE",
		X"B6",X"6D",X"55",X"15",X"22",X"04",X"41",X"20",X"08",X"11",X"49",X"92",X"24",X"A5",X"52",X"95",
		X"AA",X"B5",X"DB",X"EE",X"EE",X"EE",X"ED",X"DD",X"BD",X"DD",X"ED",X"AE",X"AD",X"B5",X"8A",X"48",
		X"20",X"40",X"00",X"41",X"10",X"11",X"12",X"49",X"A5",X"94",X"AA",X"AA",X"D5",X"ED",X"F6",X"BD",
		X"F7",X"BE",X"F7",X"7B",X"77",X"77",X"EF",X"B6",X"B5",X"55",X"55",X"10",X"41",X"10",X"40",X"10",
		X"42",X"44",X"44",X"12",X"49",X"52",X"2A",X"55",X"D5",X"DA",X"DD",X"DD",X"DB",X"F7",X"EE",X"BB",
		X"EF",X"7E",X"ED",X"75",X"5D",X"55",X"12",X"22",X"08",X"10",X"08",X"22",X"44",X"14",X"49",X"92",
		X"52",X"AA",X"54",X"D5",X"BA",X"DD",X"DE",X"7D",X"EF",X"FD",X"DD",X"BB",X"FB",X"6E",X"BB",X"AE",
		X"5A",X"0A",X"09",X"84",X"00",X"02",X"21",X"22",X"12",X"91",X"24",X"95",X"24",X"55",X"55",X"6B",
		X"BD",X"B7",X"7B",X"F7",X"DE",X"FB",X"DE",X"BD",X"FB",X"EA",X"AE",X"55",X"05",X"49",X"20",X"02",
		X"20",X"84",X"88",X"48",X"24",X"49",X"4A",X"AA",X"52",X"55",X"6D",X"B7",X"77",X"EF",X"DE",X"BB",
		X"EF",X"DB",X"7E",X"DF",X"D6",X"B7",X"5A",X"25",X"90",X"10",X"02",X"40",X"04",X"09",X"11",X"49",
		X"92",X"44",X"A5",X"52",X"55",X"D5",X"6E",X"7B",X"BB",X"6F",X"DF",X"77",X"BF",X"BB",X"BF",X"6D",
		X"BB",X"AD",X"2A",X"22",X"01",X"24",X"00",X"09",X"48",X"08",X"29",X"91",X"92",X"54",X"52",X"55",
		X"D5",X"BA",X"DD",X"ED",X"DE",X"7B",X"EF",X"7D",X"FB",X"EE",X"B7",X"DA",X"AB",X"AA",X"20",X"12",
		X"40",X"04",X"44",X"10",X"12",X"91",X"24",X"92",X"92",X"2A",X"95",X"AD",X"76",X"BB",X"FB",X"EE",
		X"BE",X"77",X"7F",X"77",X"EF",X"6E",X"AB",X"B6",X"4A",X"42",X"40",X"40",X"40",X"80",X"88",X"10",
		X"89",X"28",X"25",X"A9",X"4A",X"B5",X"AA",X"BD",X"DD",X"77",X"F7",X"7B",X"EF",X"DD",X"7B",X"B5",
		X"5B",X"B7",X"AA",X"55",X"22",X"41",X"10",X"01",X"42",X"40",X"22",X"24",X"89",X"54",X"92",X"AA",
		X"54",X"55",X"BB",X"DD",X"DD",X"BD",X"F7",X"EE",X"EE",X"6E",X"DB",X"DA",X"B6",X"55",X"55",X"55",
		X"10",X"84",X"04",X"40",X"08",X"21",X"44",X"2A",X"29",X"A5",X"AA",X"AA",X"6A",X"DD",X"ED",X"F6",
		X"BE",X"77",X"B7",X"DD",X"AD",X"6D",X"57",X"D5",X"B6",X"4A",X"55",X"9B",X"00",X"24",X"04",X"44",
		X"80",X"88",X"48",X"4A",X"51",X"95",X"54",X"AD",X"6A",X"DD",X"76",X"77",X"DF",X"DD",X"B6",X"B5",
		X"5B",X"D5",X"56",X"B5",X"5B",X"D5",X"56",X"55",X"01",X"A4",X"40",X"08",X"04",X"25",X"11",X"A5",
		X"A4",X"2A",X"55",X"AB",X"D5",X"ED",X"F6",X"76",X"EB",X"6E",X"B5",X"AD",X"D6",X"D5",X"D5",X"BA",
		X"AD",X"EA",X"AD",X"4A",X"80",X"2A",X"01",X"11",X"22",X"09",X"91",X"2A",X"49",X"95",X"AA",X"6A",
		X"D5",X"DB",X"DA",X"56",X"DB",X"AA",X"B5",X"AA",X"B5",X"76",X"2F",X"FD",X"AF",X"F4",X"D6",X"6E",
		X"09",X"29",X"22",X"12",X"21",X"92",X"44",X"52",X"92",X"B4",X"24",X"55",X"55",X"55",X"55",X"ED",
		X"A2",X"5A",X"A9",X"AA",X"EA",X"DB",X"B6",X"F7",X"BB",X"ED",X"BE",X"6B",X"95",X"22",X"25",X"90",
		X"22",X"48",X"22",X"29",X"45",X"AA",X"2A",X"55",X"55",X"55",X"25",X"55",X"95",X"AA",X"A8",X"52",
		X"5D",X"FD",X"DD",X"D6",X"FE",X"AB",X"BE",X"AB",X"AD",X"54",X"45",X"24",X"42",X"24",X"11",X"52",
		X"4A",X"92",X"AA",X"94",X"52",X"55",X"4A",X"4A",X"AA",X"4A",X"29",X"A5",X"56",X"DB",X"DF",X"BB",
		X"FE",X"BD",X"DA",X"DB",X"6D",X"29",X"55",X"49",X"44",X"88",X"28",X"89",X"24",X"45",X"AA",X"44",
		X"A5",X"4A",X"49",X"A4",X"54",X"29",X"52",X"A9",X"DA",X"6E",X"7F",X"EF",X"DA",X"FF",X"AA",X"FB",
		X"AE",X"AA",X"6A",X"55",X"48",X"52",X"44",X"94",X"24",X"92",X"54",X"09",X"A9",X"52",X"2A",X"89",
		X"AA",X"4A",X"55",X"AA",X"BA",X"AA",X"DF",X"F5",X"5D",X"FF",X"AB",X"7A",X"AF",X"AA",X"AA",X"2A",
		X"A2",X"84",X"48",X"22",X"89",X"88",X"14",X"A5",X"44",X"AA",X"AA",X"54",X"AA",X"AA",X"AA",X"AA",
		X"75",X"6B",X"F7",X"F7",X"B6",X"FB",X"BF",X"AA",X"FB",X"AA",X"AA",X"2A",X"52",X"22",X"24",X"11",
		X"42",X"52",X"84",X"A4",X"4A",X"54",X"AA",X"AA",X"4A",X"B5",X"AA",X"5A",X"D5",X"6D",X"BB",X"DD",
		X"DF",X"FA",X"DE",X"F6",X"DA",X"ED",X"4A",X"55",X"15",X"92",X"20",X"22",X"42",X"42",X"22",X"A9",
		X"28",X"A9",X"54",X"55",X"55",X"B5",X"AA",X"5B",X"BB",X"55",X"F7",X"F6",X"76",X"DB",X"BB",X"6F",
		X"AB",X"B7",X"55",X"A5",X"A2",X"04",X"81",X"44",X"08",X"11",X"49",X"24",X"49",X"AA",X"94",X"54",
		X"55",X"AD",X"AA",X"B7",X"D5",X"B6",X"DB",X"DD",X"BA",X"DF",X"D5",X"FD",X"D5",X"DA",X"B5",X"55",
		X"49",X"11",X"88",X"22",X"10",X"24",X"89",X"48",X"4A",X"4A",X"95",X"AA",X"AA",X"6A",X"6F",X"B5",
		X"DB",X"76",X"AF",X"D5",X"BB",X"75",X"57",X"DB",X"77",X"55",X"DD",X"AA",X"50",X"24",X"11",X"08",
		X"22",X"44",X"88",X"24",X"49",X"4A",X"2A",X"55",X"B5",X"75",X"DB",X"BB",X"6D",X"AF",X"DB",X"B6",
		X"ED",X"B6",X"6D",X"B7",X"5B",X"B7",X"D5",X"B6",X"12",X"12",X"01",X"42",X"20",X"84",X"48",X"24",
		X"49",X"52",X"29",X"A5",X"6A",X"55",X"F5",X"6D",X"77",X"DB",X"EE",X"AE",X"B6",X"DB",X"5A",X"57",
		X"77",X"AB",X"D6",X"AA",X"55",X"40",X"11",X"08",X"41",X"88",X"08",X"89",X"A4",X"A4",X"94",X"52",
		X"55",X"6D",X"B7",X"DD",X"DD",X"BB",X"DD",X"6D",X"B7",X"5B",X"6B",X"AB",X"BD",X"55",X"BB",X"AA",
		X"AA",X"12",X"41",X"20",X"42",X"20",X"84",X"88",X"44",X"52",X"52",X"AA",X"AA",X"AA",X"BD",X"6D",
		X"77",X"77",X"77",X"BB",X"DB",X"76",X"B7",X"D5",X"76",X"AB",X"56",X"D5",X"56",X"48",X"12",X"40",
		X"04",X"41",X"08",X"11",X"49",X"92",X"54",X"4A",X"55",X"D5",X"5A",X"BD",X"DD",X"7D",X"BB",X"BB",
		X"DD",X"B6",X"BB",X"55",X"B5",X"5D",X"55",X"55",X"A9",X"24",X"41",X"44",X"20",X"88",X"10",X"22",
		X"22",X"52",X"52",X"52",X"55",X"55",X"AB",X"BD",X"BB",X"7D",X"77",X"77",X"DB",X"DD",X"6D",X"6D",
		X"5B",X"6D",X"55",X"AB",X"A2",X"52",X"84",X"10",X"09",X"42",X"04",X"21",X"22",X"12",X"29",X"29",
		X"95",X"AA",X"5A",X"D5",X"77",X"DB",X"BD",X"77",X"77",X"B7",X"BB",X"ED",X"56",X"75",X"5B",X"95",
		X"AA",X"4A",X"89",X"10",X"89",X"20",X"42",X"84",X"90",X"44",X"92",X"94",X"54",X"95",X"AA",X"B6",
		X"EE",X"76",X"EF",X"BD",X"BD",X"7B",X"BB",X"DD",X"DA",X"D6",X"B6",X"4A",X"B5",X"2A",X"42",X"89",
		X"88",X"10",X"21",X"84",X"48",X"22",X"92",X"24",X"A5",X"AA",X"AA",X"DA",X"6D",X"77",X"EF",X"DD",
		X"BD",X"7B",X"BB",X"DD",X"D5",X"DA",X"AE",X"52",X"55",X"45",X"A4",X"44",X"20",X"22",X"22",X"82",
		X"90",X"12",X"49",X"92",X"54",X"A5",X"52",X"AD",X"DD",X"76",X"EF",X"BD",X"DB",X"FD",X"6E",X"BB",
		X"DB",X"D6",X"AA",X"D5",X"56",X"89",X"52",X"24",X"44",X"44",X"84",X"10",X"91",X"24",X"49",X"4A",
		X"4A",X"55",X"AA",X"AD",X"7A",X"B7",X"7B",X"F7",X"EE",X"BD",X"77",X"DB",X"76",X"5B",X"55",X"AD",
		X"44",X"52",X"24",X"41",X"08",X"22",X"02",X"91",X"10",X"94",X"24",X"55",X"49",X"55",X"B5",X"75",
		X"DB",X"ED",X"BB",X"FB",X"BE",X"BB",X"77",X"77",X"DB",X"DA",X"56",X"55",X"95",X"24",X"49",X"04",
		X"82",X"08",X"21",X"04",X"51",X"92",X"28",X"A9",X"52",X"A5",X"5A",X"B5",X"DB",X"F6",X"DE",X"DD",
		X"BD",X"7B",X"EF",X"6E",X"77",X"6B",X"6D",X"55",X"55",X"A4",X"24",X"88",X"10",X"22",X"10",X"12",
		X"24",X"49",X"92",X"54",X"A9",X"AA",X"AA",X"BD",X"75",X"BB",X"77",X"77",X"EF",X"DD",X"BB",X"BB",
		X"6D",X"D7",X"D6",X"AA",X"AA",X"48",X"22",X"88",X"10",X"08",X"11",X"10",X"49",X"24",X"25",X"29",
		X"95",X"AA",X"5A",X"AB",X"BB",X"DB",X"DD",X"BD",X"77",X"EF",X"F6",X"EE",X"B6",X"DB",X"DA",X"56",
		X"55",X"55",X"48",X"84",X"20",X"84",X"20",X"88",X"84",X"48",X"92",X"54",X"49",X"55",X"55",X"6D",
		X"DB",X"BD",X"BB",X"BB",X"7B",X"77",X"F7",X"DD",X"BA",X"5B",X"5B",X"AB",X"55",X"25",X"49",X"04",
		X"21",X"08",X"21",X"20",X"44",X"24",X"22",X"A5",X"52",X"A5",X"AA",X"D6",X"BA",X"ED",X"DD",X"ED",
		X"BD",X"BB",X"77",X"7B",X"77",X"DB",X"76",X"55",X"5B",X"55",X"8A",X"24",X"82",X"10",X"41",X"88",
		X"40",X"44",X"42",X"49",X"29",X"55",X"55",X"B5",X"BA",X"DD",X"EE",X"EE",X"F6",X"DD",X"DE",X"BD",
		X"B5",X"BD",X"55",X"DB",X"AA",X"54",X"51",X"44",X"10",X"22",X"04",X"82",X"10",X"52",X"10",X"55",
		X"4A",X"AA",X"AA",X"D6",X"BA",X"DB",X"DE",X"ED",X"DE",X"7B",X"BB",X"DD",X"DE",X"B5",X"BA",X"55",
		X"B5",X"4A",X"2A",X"41",X"48",X"44",X"10",X"84",X"20",X"09",X"51",X"52",X"92",X"AA",X"AA",X"5A",
		X"B7",X"BB",X"BB",X"7B",X"6F",X"77",X"F7",X"B6",X"DD",X"6E",X"5B",X"D5",X"56",X"55",X"24",X"92",
		X"10",X"22",X"08",X"21",X"88",X"44",X"24",X"89",X"52",X"95",X"AA",X"D6",X"DE",X"76",X"F7",X"76",
		X"77",X"6F",X"B7",X"DB",X"B6",X"DD",X"D6",X"AA",X"AA",X"2A",X"22",X"11",X"22",X"42",X"20",X"22",
		X"88",X"44",X"22",X"49",X"29",X"55",X"55",X"B5",X"BB",X"DD",X"BD",X"BB",X"77",X"F7",X"B6",X"BB",
		X"B5",X"6D",X"5B",X"55",X"55",X"15",X"91",X"88",X"44",X"08",X"22",X"22",X"22",X"24",X"49",X"92",
		X"54",X"AA",X"AA",X"B6",X"DB",X"BB",X"7B",X"F7",X"DD",X"DD",X"6D",X"6F",X"6B",X"DB",X"B5",X"AA",
		X"AA",X"8A",X"14",X"49",X"44",X"10",X"22",X"22",X"22",X"12",X"29",X"49",X"4A",X"A9",X"AA",X"5A",
		X"BB",X"DD",X"BD",X"7B",X"B7",X"BB",X"DB",X"6E",X"B7",X"55",X"DB",X"AA",X"94",X"54",X"44",X"24",
		X"44",X"22",X"08",X"09",X"11",X"49",X"22",X"49",X"25",X"A9",X"AA",X"DA",X"DB",X"76",X"F7",X"DD",
		X"DD",X"BD",X"BB",X"ED",X"B6",X"AD",X"B5",X"55",X"55",X"55",X"24",X"91",X"88",X"88",X"84",X"48",
		X"88",X"48",X"22",X"49",X"49",X"A5",X"AA",X"56",X"AD",X"EF",X"6E",X"B7",X"EF",X"6E",X"77",X"BB",
		X"DD",X"B6",X"5A",X"6D",X"55",X"51",X"4A",X"44",X"24",X"22",X"44",X"12",X"22",X"12",X"49",X"92",
		X"A4",X"A4",X"AA",X"AA",X"6A",X"EF",X"6E",X"7B",X"77",X"B7",X"BB",X"BB",X"5D",X"DB",X"AD",X"55",
		X"AD",X"55",X"21",X"A9",X"48",X"22",X"42",X"12",X"11",X"49",X"24",X"89",X"A4",X"54",X"4A",X"55",
		X"55",X"DB",X"BB",X"DB",X"DE",X"BB",X"DD",X"DE",X"6D",X"DB",X"76",X"AB",X"6A",X"AB",X"8A",X"22",
		X"49",X"24",X"84",X"24",X"22",X"92",X"48",X"14",X"49",X"4A",X"A5",X"AA",X"AA",X"F5",X"76",X"D7",
		X"ED",X"DE",X"76",X"77",X"DB",X"ED",X"B6",X"5B",X"55",X"B5",X"56",X"91",X"94",X"24",X"11",X"11",
		X"22",X"11",X"92",X"24",X"92",X"24",X"A9",X"54",X"AA",X"55",X"55",X"DF",X"6E",X"BB",X"DD",X"DB",
		X"6D",X"77",X"DB",X"B6",X"B6",X"AA",X"D6",X"0A",X"95",X"48",X"52",X"44",X"88",X"44",X"22",X"92",
		X"14",X"49",X"4A",X"A5",X"54",X"AA",X"6A",X"5B",X"6F",X"B7",X"BD",X"DD",X"ED",X"B6",X"BB",X"5B",
		X"77",X"B5",X"6A",X"B5",X"AA",X"8A",X"54",X"22",X"49",X"44",X"44",X"48",X"12",X"91",X"48",X"52",
		X"92",X"AA",X"52",X"D5",X"AA",X"7D",X"BB",X"DD",X"6E",X"DB",X"6E",X"DB",X"75",X"DB",X"B6",X"B6",
		X"B6",X"AA",X"4A",X"A9",X"24",X"91",X"90",X"48",X"90",X"24",X"12",X"49",X"92",X"94",X"AA",X"AA",
		X"AA",X"DA",X"DE",X"DA",X"76",X"77",X"ED",X"76",X"DB",X"B6",X"5B",X"B5",X"AD",X"55",X"15",X"55",
		X"25",X"89",X"88",X"08",X"11",X"11",X"92",X"44",X"92",X"54",X"A5",X"AA",X"AA",X"B5",X"EA",X"ED",
		X"D6",X"DD",X"6E",X"DB",X"76",X"DB",X"6E",X"DB",X"BA",X"6D",X"95",X"AA",X"A4",X"12",X"92",X"44",
		X"10",X"11",X"91",X"48",X"12",X"49",X"AA",X"52",X"55",X"55",X"DB",X"6B",X"77",X"DB",X"6E",X"B7",
		X"DD",X"6D",X"BB",X"AD",X"6D",X"6B",X"AD",X"AA",X"4A",X"29",X"49",X"44",X"08",X"11",X"12",X"89",
		X"48",X"24",X"95",X"A4",X"AA",X"54",X"55",X"6D",X"BD",X"DD",X"76",X"DB",X"DD",X"B6",X"BB",X"6D",
		X"AD",X"DD",X"5A",X"55",X"55",X"A5",X"24",X"11",X"49",X"88",X"10",X"51",X"44",X"24",X"25",X"49",
		X"A5",X"54",X"B5",X"AA",X"F5",X"6D",X"DB",X"EE",X"76",X"DB",X"DD",X"DD",X"DA",X"B6",X"6D",X"55",
		X"6B",X"55",X"95",X"24",X"49",X"88",X"88",X"88",X"44",X"84",X"52",X"92",X"52",X"4A",X"55",X"55",
		X"55",X"5B",X"6F",X"DB",X"DD",X"6E",X"B7",X"DB",X"76",X"5B",X"DD",X"B6",X"6A",X"55",X"95",X"24",
		X"25",X"24",X"11",X"12",X"12",X"11",X"91",X"24",X"49",X"4A",X"A5",X"AA",X"54",X"6B",X"D5",X"DE",
		X"EE",X"5E",X"DB",X"ED",X"B6",X"DB",X"DA",X"B6",X"AD",X"AD",X"AA",X"AA",X"A4",X"92",X"88",X"24",
		X"48",X"44",X"44",X"12",X"91",X"24",X"95",X"92",X"AA",X"AA",X"5A",X"7B",X"DB",X"76",X"77",X"B7",
		X"6D",X"77",X"BB",X"B5",X"6D",X"5B",X"AD",X"56",X"55",X"49",X"12",X"49",X"22",X"22",X"22",X"12",
		X"11",X"49",X"52",X"52",X"2A",X"55",X"55",X"55",X"5B",X"7D",X"BB",X"DD",X"ED",X"B6",X"DD",X"5D",
		X"DB",X"DA",X"B6",X"55",X"6B",X"55",X"25",X"49",X"24",X"22",X"22",X"22",X"12",X"91",X"24",X"25",
		X"49",X"55",X"4A",X"D5",X"AA",X"B5",X"5E",X"B7",X"B5",X"DB",X"DD",X"76",X"BB",X"6D",X"B7",X"6D",
		X"AD",X"B5",X"AA",X"22",X"95",X"44",X"44",X"42",X"22",X"22",X"11",X"25",X"49",X"29",X"A5",X"54",
		X"AA",X"AA",X"AA",X"ED",X"B5",X"DD",X"6D",X"B7",X"ED",X"6E",X"DB",X"B6",X"ED",X"B6",X"B5",X"AA",
		X"4A",X"92",X"48",X"48",X"22",X"22",X"49",X"92",X"28",X"25",X"A9",X"54",X"A5",X"AA",X"6A",X"AD",
		X"BE",X"6D",X"ED",X"76",X"77",X"DB",X"6E",X"6D",X"57",X"6B",X"AB",X"AA",X"52",X"52",X"12",X"91",
		X"44",X"44",X"24",X"49",X"24",X"49",X"49",X"A5",X"52",X"55",X"55",X"75",X"D5",X"B7",X"6D",X"BB",
		X"6D",X"77",X"BB",X"6D",X"6D",X"5B",X"B5",X"5A",X"55",X"25",X"15",X"89",X"48",X"12",X"11",X"89",
		X"48",X"52",X"92",X"94",X"94",X"AA",X"54",X"55",X"D5",X"DA",X"7A",X"B7",X"6D",X"DD",X"6E",X"B7",
		X"6D",X"B5",X"6B",X"55",X"AB",X"54",X"29",X"25",X"91",X"24",X"11",X"49",X"92",X"A4",X"24",X"95",
		X"2A",X"A9",X"AA",X"AA",X"5A",X"DB",X"FA",X"6E",X"DB",X"B6",X"6D",X"BB",X"B5",X"B6",X"B5",X"B6",
		X"56",X"29",X"A5",X"94",X"24",X"48",X"92",X"48",X"92",X"48",X"49",X"52",X"4A",X"2A",X"55",X"55",
		X"D5",X"DA",X"6A",X"F5",X"BB",X"B6",X"6E",X"6D",X"DB",X"B6",X"56",X"5B",X"AB",X"A4",X"2A",X"A5",
		X"24",X"89",X"88",X"94",X"48",X"92",X"44",X"52",X"49",X"2A",X"A5",X"AA",X"AA",X"D6",X"AA",X"B6",
		X"6F",X"7B",X"DB",X"B6",X"B5",X"6D",X"B7",X"B6",X"D6",X"6A",X"55",X"A9",X"A4",X"54",X"22",X"52",
		X"44",X"92",X"24",X"49",X"92",X"52",X"52",X"55",X"55",X"55",X"5B",X"5B",X"F5",X"5B",X"DB",X"B6",
		X"6D",X"DB",X"5A",X"B7",X"D5",X"5A",X"5B",X"A5",X"54",X"4A",X"55",X"09",X"91",X"24",X"91",X"24",
		X"49",X"4A",X"A5",X"24",X"55",X"55",X"B5",X"56",X"5B",X"FB",X"6E",X"6B",X"DB",X"6D",X"6D",X"6D",
		X"5D",X"5B",X"B5",X"5A",X"4A",X"A5",X"94",X"24",X"11",X"91",X"24",X"91",X"24",X"89",X"54",X"92",
		X"54",X"A9",X"AA",X"6A",X"AB",X"56",X"B5",X"6F",X"DB",X"76",X"DB",X"B6",X"5B",X"DB",X"B6",X"DA",
		X"5A",X"2B",X"55",X"52",X"29",X"09",X"91",X"48",X"92",X"24",X"92",X"24",X"49",X"29",X"25",X"95",
		X"AA",X"AA",X"D6",X"6A",X"6D",X"BF",X"B5",X"75",X"6D",X"5B",X"DB",X"6D",X"5B",X"6B",X"B5",X"6A",
		X"54",X"25",X"A5",X"14",X"49",X"24",X"25",X"4A",X"2A",X"4A",X"29",X"A9",X"AA",X"AA",X"5A",X"AB",
		X"AA",X"56",X"EB",X"B6",X"55",X"A9",X"2A",X"2D",X"4B",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"66",X"AB",X"A4",X"AA",X"4A",X"A9",X"CA",X"CA",X"54",X"99",X"B1",X"AA",X"CA",X"99",
		X"C9",X"9A",X"A9",X"B2",X"32",X"D9",X"A4",X"AA",X"92",X"59",X"B5",X"AA",X"66",X"5A",X"69",X"51",
		X"AB",X"A8",X"68",X"4A",X"52",X"A5",X"96",X"17",X"6A",X"B5",X"96",X"45",X"5A",X"DA",X"92",X"6A",
		X"35",X"69",X"B5",X"CA",X"AA",X"B4",X"B4",X"96",X"AE",X"B2",X"55",X"25",X"4A",X"5D",X"A9",X"D4",
		X"56",X"69",X"AD",X"5E",X"B7",X"A4",X"5F",X"57",X"EB",X"BE",X"AA",X"AA",X"5A",X"D5",X"A9",X"28",
		X"D7",X"D5",X"2B",X"0A",X"25",X"49",X"28",X"84",X"16",X"6A",X"FD",X"9F",X"08",X"00",X"80",X"6A",
		X"81",X"97",X"FF",X"FF",X"01",X"00",X"00",X"FE",X"D7",X"01",X"BC",X"FF",X"0F",X"00",X"00",X"F8",
		X"FF",X"07",X"00",X"FE",X"FF",X"03",X"00",X"F8",X"FF",X"07",X"00",X"FC",X"FF",X"0F",X"00",X"E0",
		X"FF",X"07",X"00",X"FC",X"FF",X"03",X"00",X"F8",X"FF",X"01",X"00",X"FF",X"7F",X"00",X"00",X"FF",
		X"3F",X"00",X"C0",X"FF",X"0F",X"00",X"E0",X"FF",X"03",X"00",X"F8",X"FF",X"01",X"00",X"FE",X"3F",
		X"00",X"80",X"FF",X"0F",X"00",X"E0",X"FF",X"03",X"00",X"FC",X"FF",X"00",X"00",X"FF",X"1F",X"00",
		X"C0",X"FF",X"07",X"00",X"F8",X"FF",X"00",X"00",X"FE",X"3F",X"00",X"E0",X"FF",X"07",X"00",X"F8",
		X"FF",X"08",X"80",X"FF",X"1F",X"00",X"E0",X"FF",X"33",X"00",X"FE",X"7F",X"00",X"C0",X"FF",X"37",
		X"00",X"FC",X"FF",X"00",X"C0",X"FF",X"77",X"00",X"F0",X"FF",X"01",X"C0",X"FF",X"7F",X"00",X"E0",
		X"FF",X"01",X"E0",X"FF",X"3D",X"00",X"F8",X"7F",X"00",X"F0",X"7F",X"0F",X"00",X"FC",X"1F",X"00",
		X"FC",X"DF",X"03",X"80",X"DF",X"C7",X"00",X"FF",X"7B",X"00",X"E0",X"FF",X"19",X"F0",X"3F",X"0F",
		X"00",X"FE",X"8F",X"00",X"FF",X"77",X"00",X"F0",X"FF",X"08",X"E0",X"FF",X"07",X"00",X"FE",X"FF",
		X"00",X"FE",X"77",X"00",X"C0",X"FD",X"1F",X"F0",X"9F",X"03",X"00",X"CC",X"E7",X"C0",X"FF",X"1E",
		X"00",X"60",X"EF",X"01",X"FE",X"F7",X"00",X"00",X"7B",X"1E",X"F8",X"DF",X"03",X"00",X"10",X"3D",
		X"F0",X"7F",X"07",X"80",X"60",X"70",X"E0",X"7F",X"0F",X"00",X"82",X"E3",X"01",X"F9",X"3F",X"04",
		X"00",X"F1",X"0D",X"FE",X"3F",X"0C",X"02",X"E0",X"0B",X"FF",X"3F",X"00",X"0E",X"C3",X"18",X"FF",
		X"3F",X"00",X"06",X"E3",X"9A",X"FF",X"1F",X"00",X"43",X"70",X"1C",X"FF",X"0F",X"80",X"C0",X"F8",
		X"58",X"FF",X"07",X"20",X"00",X"7E",X"FF",X"FF",X"00",X"38",X"04",X"C7",X"FF",X"7F",X"00",X"82",
		X"E0",X"F6",X"FF",X"0F",X"C0",X"20",X"38",X"FD",X"FF",X"03",X"30",X"00",X"AF",X"FF",X"3F",X"00",
		X"86",X"E0",X"6D",X"FF",X"0F",X"C0",X"20",X"B8",X"FF",X"FF",X"00",X"94",X"02",X"E9",X"FF",X"3F",
		X"02",X"44",X"70",X"BC",X"FF",X"1F",X"08",X"00",X"DA",X"FB",X"FF",X"41",X"0A",X"00",X"AD",X"FF",
		X"7F",X"80",X"04",X"A8",X"FA",X"FF",X"07",X"42",X"80",X"AA",X"FB",X"FF",X"02",X"02",X"90",X"F5",
		X"FF",X"1F",X"20",X"04",X"B2",X"FE",X"FF",X"0B",X"04",X"80",X"EC",X"FE",X"FF",X"10",X"04",X"50",
		X"ED",X"FF",X"3F",X"20",X"02",X"D8",X"FE",X"FF",X"05",X"21",X"40",X"D5",X"FF",X"7F",X"01",X"11",
		X"90",X"F6",X"FF",X"5F",X"20",X"04",X"A8",X"ED",X"FF",X"2F",X"08",X"01",X"D2",X"FE",X"FF",X"8B",
		X"08",X"04",X"65",X"F7",X"FF",X"96",X"22",X"40",X"D4",X"FE",X"7D",X"2B",X"55",X"02",X"48",X"AB",
		X"DA",X"BB",X"B6",X"4A",X"A2",X"2A",X"45",X"69",X"5F",X"A5",X"F6",X"5A",X"AA",X"5A",X"D5",X"B9",
		X"40",X"DC",X"57",X"77",X"AF",X"AA",X"95",X"48",X"AB",X"F5",X"5E",X"AD",X"6A",X"6B",X"AB",X"45",
		X"E9",X"EB",X"42",X"E5",X"B7",X"52",X"54",X"75",X"1E",X"9B",X"2B",X"2A",X"AD",X"51",X"F5",X"AB",
		X"A2",X"54",X"95",X"A2",X"BA",X"57",X"15",X"95",X"AA",X"94",X"D6",X"B5",X"15",X"A5",X"BA",X"AE",
		X"4A",X"69",X"5D",X"AA",X"EA",X"FA",X"AE",X"CA",X"E9",X"BA",X"AA",X"F5",X"DA",X"AA",X"6A",X"D5",
		X"DA",X"F6",X"6A",X"55",X"55",X"35",X"AA",X"5E",X"6F",X"55",X"28",X"A5",X"52",X"55",X"5F",X"D7",
		X"2A",X"94",X"4A",X"A9",X"54",X"DB",X"A5",X"28",X"2A",X"4B",X"A9",X"5A",X"AB",X"52",X"AA",X"4E",
		X"AB",X"52",X"52",X"55",X"63",X"A9",X"5E",X"97",X"B2",X"AA",X"4E",X"55",X"75",X"2D",X"D1",X"7A",
		X"5B",X"95",X"52",X"55",X"AB",X"EA",X"BB",X"5A",X"45",X"A9",X"AA",X"D6",X"AA",X"2A",X"8A",X"AA",
		X"54",X"D5",X"D6",X"51",X"2A",X"55",X"AB",X"2A",X"2A",X"A5",X"A2",X"54",X"57",X"A5",X"5A",X"95",
		X"52",X"75",X"55",X"55",X"D1",X"54",X"55",X"E3",X"A8",X"56",X"AB",X"52",X"B5",X"56",X"65",X"55",
		X"95",X"56",X"51",X"55",X"AB",X"AA",X"5A",X"55",X"51",X"15",X"AD",X"EB",X"5D",X"AD",X"44",X"A9",
		X"54",X"56",X"EB",X"29",X"0A",X"C7",X"71",X"CE",X"73",X"CE",X"E3",X"70",X"CE",X"79",X"1C",X"3C",
		X"73",X"78",X"7A",X"9E",X"17",X"8E",X"38",X"8E",X"E1",X"9D",X"F3",X"18",X"E6",X"38",X"C6",X"39",
		X"8E",X"83",X"54",X"20",X"DE",X"61",X"5E",X"86",X"A9",X"32",X"B3",X"2C",X"E3",X"38",X"E6",X"71",
		X"8E",X"66",X"9C",X"52",X"8E",X"63",X"8C",X"69",X"1C",X"B7",X"99",X"23",X"CC",X"CC",X"75",X"6C",
		X"57",X"B3",X"D8",X"A8",X"56",X"D6",X"36",X"CE",X"B5",X"B8",X"EF",X"EF",X"3C",X"43",X"08",X"82",
		X"52",X"46",X"E7",X"F1",X"DE",X"FF",X"9E",X"93",X"00",X"00",X"81",X"52",X"9B",X"1D",X"EF",X"FA",
		X"FE",X"DF",X"4A",X"00",X"00",X"10",X"4E",X"DB",X"6E",X"DB",X"EE",X"FF",X"BF",X"2D",X"00",X"00",
		X"80",X"E9",X"6E",X"CF",X"B5",X"F6",X"7F",X"FF",X"53",X"00",X"00",X"00",X"E9",X"DE",X"E7",X"69",
		X"AD",X"FF",X"FF",X"4D",X"00",X"00",X"00",X"70",X"EF",X"EF",X"AA",X"2A",X"EF",X"FF",X"6F",X"01",
		X"00",X"00",X"C0",X"FA",X"FB",X"56",X"A5",X"EA",X"FF",X"7F",X"0F",X"00",X"00",X"00",X"7A",X"FF",
		X"9F",X"2D",X"8C",X"FD",X"FF",X"E7",X"01",X"00",X"00",X"C0",X"F7",X"FF",X"E3",X"42",X"D1",X"FF",
		X"EF",X"73",X"00",X"00",X"00",X"E8",X"FF",X"FF",X"55",X"41",X"E2",X"FB",X"FF",X"E3",X"00",X"00",
		X"00",X"F0",X"FF",X"FF",X"57",X"01",X"A1",X"FF",X"FF",X"8F",X"03",X"00",X"00",X"8C",X"FF",X"FF",
		X"3F",X"06",X"00",X"EF",X"FF",X"FF",X"31",X"00",X"00",X"C0",X"FF",X"FF",X"57",X"01",X"00",X"80",
		X"FF",X"FF",X"EF",X"01",X"00",X"00",X"E0",X"FF",X"7F",X"03",X"00",X"00",X"EA",X"FF",X"FF",X"3F",
		X"07",X"00",X"00",X"FC",X"FF",X"7F",X"00",X"00",X"80",X"FD",X"FF",X"FF",X"3F",X"18",X"00",X"00",
		X"FC",X"FF",X"FF",X"01",X"00",X"80",X"FE",X"FF",X"DF",X"FF",X"0F",X"0F",X"04",X"00",X"FD",X"FF",
		X"79",X"00",X"00",X"C0",X"EF",X"DF",X"A7",X"FD",X"1F",X"0F",X"00",X"00",X"FE",X"FF",X"73",X"00",
		X"00",X"F0",X"7F",X"3F",X"0E",X"FE",X"7F",X"3E",X"00",X"00",X"E0",X"FF",X"1F",X"02",X"00",X"40",
		X"FD",X"DF",X"05",X"95",X"FF",X"BF",X"07",X"00",X"00",X"FD",X"FF",X"03",X"00",X"00",X"F8",X"FF",
		X"03",X"05",X"DC",X"FF",X"9F",X"03",X"00",X"C0",X"FF",X"FF",X"03",X"00",X"60",X"F3",X"F7",X"01",
		X"10",X"FC",X"FF",X"3F",X"04",X"00",X"80",X"FF",X"FF",X"05",X"00",X"00",X"FF",X"7F",X"09",X"00",
		X"D6",X"FF",X"FF",X"03",X"00",X"00",X"FD",X"FF",X"0F",X"00",X"00",X"FD",X"FF",X"1F",X"00",X"00",
		X"FE",X"FF",X"FF",X"03",X"00",X"80",X"FE",X"FF",X"17",X"00",X"80",X"FE",X"FF",X"0B",X"00",X"00",
		X"FC",X"FF",X"FF",X"7F",X"00",X"00",X"D0",X"FD",X"5F",X"04",X"00",X"A0",X"FF",X"5F",X"01",X"00",
		X"10",X"FD",X"FF",X"EF",X"FD",X"03",X"00",X"C0",X"EB",X"FF",X"42",X"00",X"40",X"FB",X"FF",X"25",
		X"00",X"00",X"BC",X"FF",X"7F",X"EF",X"1B",X"00",X"00",X"FE",X"FF",X"0A",X"00",X"40",X"FF",X"FF",
		X"85",X"00",X"00",X"D0",X"FF",X"7F",X"E5",X"FF",X"01",X"00",X"40",X"F7",X"FF",X"09",X"00",X"D0",
		X"FE",X"77",X"01",X"00",X"E0",X"7F",X"FF",X"4A",X"FF",X"FE",X"00",X"00",X"E0",X"FD",X"7D",X"08",
		X"00",X"DA",X"5F",X"95",X"80",X"C4",X"DC",X"EE",X"DD",X"FE",X"FF",X"07",X"00",X"00",X"FF",X"FF",
		X"01",X"00",X"A0",X"3F",X"FF",X"02",X"01",X"C8",X"FB",X"F7",X"FF",X"FF",X"07",X"00",X"00",X"FF",
		X"7F",X"01",X"00",X"40",X"FD",X"BF",X"0A",X"00",X"D0",X"FD",X"FF",X"EF",X"FF",X"05",X"00",X"80",
		X"FE",X"D7",X"02",X"00",X"A8",X"FE",X"77",X"45",X"00",X"E8",X"DF",X"FF",X"FF",X"BF",X"01",X"00",
		X"60",X"7F",X"AB",X"20",X"40",X"6A",X"DF",X"5B",X"02",X"50",X"ED",X"FF",X"FF",X"FF",X"02",X"00",
		X"20",X"BD",X"2D",X"22",X"04",X"AB",X"5D",X"57",X"41",X"A0",X"F6",X"FF",X"FF",X"BF",X"A5",X"00",
		X"80",X"48",X"75",X"08",X"49",X"D2",X"AE",X"D6",X"0A",X"44",X"6B",X"F7",X"FF",X"FF",X"AF",X"08",
		X"10",X"80",X"92",X"92",X"42",X"A9",X"AA",X"F5",X"5A",X"40",X"58",X"F7",X"FD",X"FF",X"6F",X"AB",
		X"04",X"01",X"08",X"22",X"4A",X"8B",X"B2",X"D5",X"EA",X"8A",X"40",X"71",X"F9",X"FF",X"7F",X"5E",
		X"D7",X"2A",X"01",X"20",X"10",X"AA",X"AA",X"D6",X"52",X"75",X"05",X"54",X"55",X"FD",X"FF",X"FF",
		X"AF",X"B5",X"08",X"00",X"01",X"A0",X"52",X"69",X"AB",X"D2",X"2A",X"48",X"55",X"F5",X"FF",X"FF",
		X"BF",X"AB",X"14",X"02",X"02",X"81",X"50",X"D5",X"6A",X"55",X"15",X"52",X"AA",X"6E",X"FF",X"FF",
		X"7E",X"AF",X"AA",X"04",X"00",X"44",X"A0",X"D4",X"52",X"55",X"4D",X"A0",X"54",X"B5",X"FE",X"FD",
		X"EF",X"BD",X"9D",X"22",X"00",X"08",X"11",X"A5",X"55",X"A9",X"5A",X"0A",X"94",X"AA",X"DD",X"EF",
		X"FF",X"ED",X"DE",X"8A",X"42",X"01",X"44",X"22",X"D5",X"A4",X"B4",X"2A",X"A2",X"54",X"D5",X"FE",
		X"F7",X"FD",X"BD",X"DB",X"45",X"29",X"04",X"22",X"A9",X"54",X"55",X"55",X"A5",X"AA",X"5A",X"EF",
		X"7B",X"7B",X"5F",X"D7",X"52",X"20",X"12",X"08",X"48",X"A8",X"94",X"54",X"A9",X"94",X"AA",X"F6",
		X"7A",X"BD",X"BB",X"EB",X"2A",X"01",X"95",X"20",X"24",X"12",X"AA",X"52",X"52",X"AA",X"AA",X"52",
		X"FD",X"BE",X"ED",X"7E",X"AD",X"94",X"4A",X"E3",X"F1",X"54",X"A5",X"2A",X"4D",X"47",X"D5",X"9A",
		X"AA",X"55",X"45",X"75",X"61",X"B5",X"5E",X"A3",X"F4",X"A8",X"58",X"1D",X"E3",X"78",X"94",X"C6",
		X"71",X"5C",X"8E",X"E3",X"28",X"CB",X"EA",X"68",X"2E",X"54",X"CB",X"E2",X"33",X"BA",X"58",X"55",
		X"B1",X"CE",X"AA",X"73",X"A8",X"0B",X"A7",X"32",X"33",X"0C",X"17",X"1D",X"C6",X"52",X"2A",X"C3",
		X"39",X"4A",X"55",X"87",X"9D",X"E3",X"9A",X"79",X"EE",X"CC",X"B9",X"66",X"DE",X"B3",X"6E",X"CE",
		X"B9",X"6A",X"F6",X"31",X"C7",X"30",X"26",X"65",X"0C",X"50",X"42",X"62",X"31",X"0A",X"1D",X"89",
		X"6B",X"8D",X"77",X"75",X"33",X"27",X"77",X"73",X"A5",X"6A",X"1F",X"66",X"27",X"23",X"D3",X"4C",
		X"76",X"A9",X"12",X"46",X"86",X"29",X"8A",X"48",X"20",X"62",X"85",X"A8",X"73",X"77",X"7E",X"BD",
		X"EB",X"97",X"EC",X"B4",X"D5",X"82",X"02",X"00",X"64",X"C5",X"18",X"C3",X"1C",X"0C",X"FB",X"01",
		X"BE",X"9D",X"FD",X"AE",X"F1",X"7F",X"DE",X"3B",X"7F",X"DE",X"BF",X"ED",X"EB",X"F6",X"D5",X"3B",
		X"DB",X"3E",X"37",X"DD",X"EC",X"72",X"77",X"A5",X"14",X"33",X"C3",X"8C",X"22",X"0E",X"00",X"19",
		X"91",X"A0",X"4C",X"10",X"11",X"22",X"50",X"01",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"99",X"B5",X"7C",X"EE",X"FD",X"DB",X"EF",X"7E",X"FF",X"FB",X"FF",X"7D",
		X"7F",X"FF",X"FD",X"FF",X"76",X"FF",X"EF",X"EF",X"EF",X"F6",X"BB",X"DE",X"EA",X"59",X"F9",X"11",
		X"5D",X"C9",X"0D",X"E2",X"C5",X"24",X"52",X"88",X"04",X"29",X"10",X"49",X"44",X"C9",X"10",X"19",
		X"52",X"51",X"4B",X"2D",X"E9",X"8E",X"B4",X"6D",X"82",X"75",X"2F",X"BA",X"91",X"0E",X"10",X"AE",
		X"98",X"77",X"75",X"04",X"56",X"D7",X"00",X"6A",X"AD",X"FB",X"7F",X"40",X"3F",X"00",X"FC",X"8F",
		X"EC",X"32",X"26",X"93",X"8C",X"07",X"25",X"9A",X"00",X"7C",X"48",X"C5",X"03",X"75",X"51",X"31",
		X"D0",X"A8",X"E2",X"2A",X"AA",X"08",X"B8",X"20",X"02",X"C0",X"04",X"DC",X"2E",X"E1",X"4C",X"D1",
		X"6A",X"57",X"DD",X"6D",X"55",X"BB",X"DF",X"F5",X"BE",X"F6",X"BD",X"AD",X"BE",X"93",X"FF",X"5C",
		X"FD",X"F3",X"F7",X"37",X"8F",X"00",X"FC",X"FF",X"FF",X"BF",X"82",X"34",X"DD",X"7B",X"E5",X"1F",
		X"DB",X"CB",X"1F",X"F0",X"5F",X"DF",X"07",X"7B",X"A2",X"8D",X"99",X"CC",X"64",X"12",X"05",X"6C",
		X"22",X"A0",X"22",X"00",X"2A",X"00",X"C0",X"20",X"42",X"05",X"12",X"18",X"08",X"90",X"4A",X"D5",
		X"44",X"74",X"A9",X"0A",X"B7",X"71",X"8F",X"EF",X"DD",X"E7",X"5B",X"7F",X"FD",X"7F",X"FA",X"FB",
		X"5E",X"3B",X"D9",X"8F",X"62",X"92",X"2A",X"06",X"BA",X"83",X"15",X"67",X"58",X"85",X"41",X"B8",
		X"81",X"27",X"3C",X"88",X"57",X"74",X"60",X"2E",X"07",X"7F",X"8C",X"B5",X"61",X"97",X"28",X"C2",
		X"00",X"0A",X"A8",X"00",X"80",X"48",X"03",X"A9",X"88",X"59",X"11",X"BD",X"89",X"FB",X"FF",X"FF",
		X"FF",X"FF",X"FB",X"EF",X"DF",X"EF",X"7B",X"EF",X"BD",X"77",X"77",X"77",X"BB",X"DD",X"6E",X"DB",
		X"B6",X"AD",X"F5",X"FF",X"FF",X"F7",X"2F",X"44",X"29",X"10",X"08",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"44",X"44",X"24",X"49",X"52",X"52",X"A9",X"AA",
		X"AA",X"D6",X"B6",X"ED",X"EE",X"EE",X"7D",X"EF",X"BD",X"F7",X"5D",X"F9",X"C4",X"B4",X"E9",X"C7",
		X"FF",X"EE",X"ED",X"7E",X"EF",X"FE",X"7F",X"BF",X"FD",X"AD",X"DB",X"FF",X"DF",X"EF",X"B6",X"37",
		X"5F",X"DA",X"B3",X"3E",X"6D",X"B6",X"29",X"D9",X"16",X"68",X"FF",X"6D",X"FB",X"0F",X"BD",X"65",
		X"68",X"42",X"04",X"08",X"00",X"00",X"00",X"00",X"BE",X"02",X"00",X"00",X"00",X"00",X"11",X"00",
		X"4C",X"00",X"A8",X"02",X"C0",X"26",X"40",X"15",X"54",X"C9",X"54",X"1D",X"DD",X"5E",X"D5",X"DD",
		X"BB",X"7F",X"BF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"BF",X"7F",X"DF",X"BB",X"77",
		X"77",X"BB",X"6D",X"B7",X"6D",X"AD",X"B5",X"56",X"AD",X"AA",X"AA",X"52",X"CA",X"6E",X"BF",X"0B",
		X"D0",X"0F",X"C8",X"50",X"1A",X"00",X"50",X"00",X"2C",X"01",X"57",X"00",X"00",X"00",X"50",X"92",
		X"02",X"F4",X"3F",X"00",X"40",X"28",X"01",X"5C",X"53",X"50",X"89",X"1E",X"42",X"7F",X"42",X"2C",
		X"97",X"60",X"BD",X"68",X"DE",X"AA",X"B2",X"17",X"68",X"6B",X"E9",X"5D",X"AD",X"F2",X"EB",X"EE",
		X"EA",X"BF",X"DD",X"77",X"FB",X"EF",X"FE",X"7B",X"FF",X"7A",X"5F",X"AF",X"FF",X"BC",X"DD",X"B6",
		X"2E",X"AD",X"AB",X"E8",X"B2",X"00",X"37",X"25",X"48",X"47",X"10",X"2A",X"48",X"16",X"84",X"41",
		X"04",X"55",X"10",X"51",X"64",X"22",X"48",X"35",X"A9",X"EE",X"6E",X"07",X"00",X"00",X"DA",X"B6",
		X"08",X"EE",X"01",X"14",X"04",X"80",X"72",X"20",X"47",X"40",X"2A",X"A0",X"14",X"CC",X"50",X"12",
		X"33",X"88",X"6E",X"52",X"9F",X"49",X"6E",X"B6",X"DD",X"AD",X"FA",X"DA",X"5D",X"75",X"7D",X"65",
		X"FE",X"3B",X"FE",X"FB",X"F2",X"F8",X"A7",X"FF",X"9F",X"EE",X"B7",X"BE",X"6F",X"C9",X"5F",X"EB",
		X"DD",X"5C",X"9F",X"AE",X"BC",X"DA",X"6A",X"31",X"F5",X"85",X"A3",X"3A",X"90",X"9C",X"CC",X"0C",
		X"A8",X"22",X"48",X"04",X"6E",X"00",X"19",X"41",X"06",X"24",X"41",X"4D",X"51",X"FC",X"FF",X"01",
		X"00",X"50",X"B7",X"EF",X"AD",X"1A",X"05",X"40",X"11",X"8A",X"E2",X"1D",X"84",X"61",X"21",X"8A",
		X"C1",X"5D",X"25",X"74",X"0B",X"E5",X"3E",X"F2",X"1D",X"9B",X"53",X"D5",X"DE",X"A8",X"FB",X"22",
		X"BD",X"CA",X"FE",X"92",X"FD",X"93",X"2B",X"AF",X"C9",X"5E",X"53",X"B7",X"55",X"FF",X"51",X"ED",
		X"DA",X"5A",X"54",X"15",X"9D",X"AD",X"5D",X"4B",X"36",X"93",X"94",X"C9",X"16",X"CA",X"16",X"26",
		X"6A",X"2E",X"22",X"CA",X"9A",X"7B",X"29",X"60",X"49",X"0D",X"FB",X"80",X"2C",X"93",X"20",X"44",
		X"00",X"20",X"15",X"E0",X"FF",X"00",X"00",X"A0",X"EE",X"5E",X"55",X"A5",X"24",X"11",X"40",X"44",
		X"DD",X"FF",X"FF",X"14",X"C7",X"30",X"BE",X"B7",X"D9",X"3C",X"EB",X"96",X"FB",X"9D",X"74",X"2F",
		X"AD",X"67",X"EB",X"5A",X"FD",X"4A",X"3B",X"95",X"F9",X"8B",X"3B",X"D7",X"DC",X"55",X"55",X"E8",
		X"36",X"5C",X"86",X"5A",X"89",X"6A",X"27",X"B9",X"48",X"16",X"C1",X"48",X"64",X"A2",X"66",X"46",
		X"A6",X"48",X"34",X"8D",X"A2",X"C1",X"D2",X"8C",X"64",X"25",X"D2",X"90",X"48",X"A1",X"0A",X"8B",
		X"6A",X"07",X"EA",X"93",X"AC",X"EF",X"E8",X"76",X"5F",X"5D",X"7F",X"FC",X"13",X"3F",X"00",X"50",
		X"EB",X"F7",X"D6",X"AA",X"10",X"09",X"89",X"88",X"22",X"15",X"28",X"66",X"9A",X"02",X"EA",X"38",
		X"0C",X"C7",X"20",X"9E",X"7B",X"CC",X"5B",X"DA",X"59",X"D6",X"BC",X"CA",X"B6",X"6B",X"CE",X"EE",
		X"4D",X"FD",X"6D",X"F6",X"73",X"FC",X"9D",X"B5",X"33",X"7F",X"DA",X"55",X"EB",X"2C",X"AB",X"79",
		X"A5",X"9F",X"A4",X"6B",X"55",X"20",X"22",X"4A",X"55",X"30",X"C9",X"A8",X"49",X"24",X"4A",X"14",
		X"25",X"D2",X"4C",X"59",X"26",X"53",X"B3",X"D2",X"A1",X"BB",X"B2",X"ED",X"06",X"E0",X"0A",X"59",
		X"26",X"21",X"19",X"24",X"B5",X"40",X"D5",X"02",X"1E",X"FF",X"38",X"00",X"00",X"D4",X"BB",X"5B",
		X"4D",X"25",X"49",X"92",X"24",X"55",X"5B",X"F7",X"BA",X"55",X"EF",X"EA",X"5C",X"0D",X"D6",X"EB",
		X"BD",X"AF",X"E3",X"BB",X"ED",X"5E",X"67",X"3D",X"D7",X"3B",X"77",X"DD",X"36",X"B3",X"F9",X"AD",
		X"3A",X"57",X"F6",X"5A",X"56",X"AF",X"B2",X"A3",X"9E",X"BA",X"E8",X"25",X"15",X"93",X"4C",X"59",
		X"E8",X"14",X"42",X"0F",X"18",X"16",X"91",X"08",X"85",X"A8",X"88",X"8C",X"4C",X"A4",X"28",X"89",
		X"2A",X"49",X"49",X"92",X"A5",X"24",X"31",X"CC",X"94",X"CA",X"6C",X"30",X"12",X"49",X"55",X"65",
		X"82",X"AE",X"44",X"E6",X"15",X"91",X"56",X"45",X"5B",X"DA",X"F8",X"5F",X"7F",X"00",X"40",X"B7",
		X"FF",X"DD",X"B6",X"B5",X"AA",X"56",X"55",X"B5",X"DD",X"F6",X"B6",X"ED",X"DA",X"6A",X"55",X"05",
		X"C0",X"CA",X"EB",X"7F",X"AB",X"22",X"2A",X"CC",X"75",X"BB",X"53",X"4C",X"13",X"B5",X"5A",X"63",
		X"57",X"D8",X"99",X"D4",X"99",X"51",X"9D",X"49",X"75",X"A1",X"99",X"1A",X"99",X"5B",X"D0",X"C3",
		X"84",X"35",X"F0",X"4C",X"8A",X"2B",X"82",X"8B",X"A5",X"C1",X"54",X"94",X"55",X"A2",X"52",X"AA",
		X"56",X"55",X"5B",X"AA",X"AA",X"EA",X"55",X"5D",X"D5",X"B6",X"DD",X"B6",X"B6",X"AA",X"DB",X"16",
		X"DD",X"66",X"F6",X"B9",X"89",X"DB",X"6A",X"C7",X"46",X"2B",X"55",X"4D",X"16",X"71",X"5F",X"DD",
		X"F5",X"0F",X"00",X"50",X"DA",X"7E",X"AD",X"55",X"95",X"A4",X"24",X"49",X"A9",X"AA",X"76",X"6D",
		X"D7",X"AA",X"2A",X"4A",X"25",X"89",X"54",X"55",X"AD",X"55",X"05",X"08",X"F4",X"75",X"DF",X"43",
		X"28",X"4D",X"F5",X"5E",X"A5",X"5A",X"45",X"75",X"67",X"5C",X"25",X"AA",X"45",X"AA",X"4A",X"D4",
		X"51",X"32",X"23",X"B2",X"A5",X"B8",X"4A",X"64",X"99",X"61",X"36",X"D1",X"66",X"B2",X"DD",X"98",
		X"D7",X"B2",X"A0",X"2B",X"E8",X"54",X"B6",X"B6",X"55",X"A5",X"AA",X"6A",X"2B",X"75",X"6D",X"75",
		X"BB",X"B6",X"56",X"55",X"B5",X"6E",X"66",X"65",X"52",X"D2",X"A6",X"CC",X"2A",X"46",X"8C",X"44",
		X"D2",X"A4",X"12",X"C9",X"94",X"8A",X"54",X"D5",X"FD",X"03",X"00",X"50",X"6A",X"DB",X"D5",X"AA",
		X"92",X"92",X"A4",X"54",X"55",X"AD",X"AB",X"6D",X"5B",X"5B",X"AD",X"AA",X"4A",X"55",X"F5",X"EE",
		X"6E",X"BB",X"ED",X"56",X"5B",X"6D",X"DB",X"ED",X"76",X"DB",X"B6",X"02",X"70",X"9D",X"EF",X"7F",
		X"C6",X"54",X"48",X"FF",X"5A",X"EB",X"28",X"52",X"2D",X"D5",X"25",X"45",X"95",X"12",X"A9",X"22",
		X"53",X"16",X"51",X"51",X"85",X"4A",X"54",X"29",X"51",X"92",X"A8",X"D8",X"28",X"45",X"85",X"8C",
		X"A4",X"52",X"91",X"2A",X"53",X"99",X"49",X"99",X"A8",X"52",X"53",X"AB",X"5A",X"DD",X"5A",X"6D",
		X"AD",X"EE",X"5A",X"77",X"55",X"5B",X"75",X"D5",X"AA",X"B5",X"AD",X"ED",X"5A",X"AB",X"5A",X"4A",
		X"55",X"EB",X"B7",X"AA",X"00",X"54",X"B5",X"F5",X"B6",X"AA",X"55",X"29",X"55",X"55",X"55",X"55",
		X"AB",X"AA",X"AA",X"AA",X"AA",X"AA",X"52",X"A4",X"52",X"55",X"B5",X"AA",X"4A",X"95",X"52",X"4A",
		X"A2",X"54",X"2A",X"55",X"52",X"55",X"25",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",
		X"20",X"AE",X"E7",X"7B",X"87",X"52",X"8A",X"F5",X"5D",X"D5",X"5A",X"42",X"B5",X"AA",X"7A",X"2D",
		X"AA",X"AA",X"A4",X"6A",X"A5",X"5A",X"55",X"55",X"A9",X"54",X"AB",X"52",X"35",X"4B",X"A9",X"54",
		X"29",X"51",X"C4",X"8C",X"95",X"52",X"8A",X"99",X"5A",X"B5",X"AA",X"4A",X"55",X"55",X"A5",X"AA",
		X"B5",X"76",X"97",X"AA",X"54",X"D5",X"EA",X"AD",X"B5",X"54",X"55",X"55",X"55",X"55",X"55",X"7D",
		X"AD",X"02",X"AA",X"AA",X"EA",X"AD",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"54",X"AA",X"AA",X"AA",X"A4",X"94",X"A4",X"54",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"49",X"4A",X"A9",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"D5",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"02",
		X"80",X"BE",X"7F",X"77",X"AB",X"AA",X"84",X"D4",X"01",X"00",X"00",X"84",X"A4",X"AA",X"ED",X"EF",
		X"FF",X"FB",X"D6",X"BF",X"BF",X"77",X"8F",X"23",X"00",X"00",X"20",X"10",X"82",X"A8",X"B6",X"7B",
		X"EF",X"BB",X"B7",X"6D",X"AB",X"75",X"97",X"84",X"88",X"48",X"4A",X"A5",X"EE",X"FF",X"FF",X"FF",
		X"EE",X"B6",X"2A",X"45",X"10",X"04",X"00",X"00",X"40",X"88",X"10",X"51",X"D5",X"B6",X"BB",X"F7",
		X"EF",X"BF",X"DF",X"77",X"DB",X"5A",X"95",X"40",X"00",X"80",X"40",X"22",X"AA",X"FB",X"FD",X"EF",
		X"F7",X"DE",X"76",X"2D",X"09",X"21",X"08",X"91",X"A4",X"54",X"D5",X"DA",X"B6",X"B6",X"B5",X"AA",
		X"2A",X"22",X"08",X"20",X"22",X"89",X"08",X"04",X"02",X"0C",X"12",X"55",X"DB",X"F7",X"F7",X"77",
		X"EF",X"FB",X"FF",X"FE",X"BE",X"AF",X"D7",X"56",X"95",X"14",X"A9",X"AA",X"B6",X"56",X"55",X"92",
		X"08",X"00",X"00",X"00",X"00",X"42",X"48",X"55",X"6B",X"EB",X"B6",X"B6",X"B5",X"B5",X"6D",X"BB",
		X"BD",X"6D",X"5D",X"AD",X"5A",X"AD",X"FB",X"FF",X"FF",X"FB",X"F7",X"6E",X"2D",X"25",X"21",X"84",
		X"20",X"04",X"08",X"00",X"40",X"20",X"AA",X"76",X"EF",X"F7",X"DD",X"5D",X"A5",X"10",X"21",X"29",
		X"55",X"55",X"AD",X"D6",X"DA",X"DA",X"76",X"A6",X"10",X"22",X"A9",X"6A",X"F5",X"FF",X"FF",X"FF",
		X"FF",X"DE",X"B6",X"52",X"82",X"40",X"40",X"00",X"10",X"40",X"10",X"92",X"94",X"6A",X"BF",X"FF",
		X"FF",X"F7",X"BD",X"B5",X"12",X"11",X"10",X"88",X"A0",X"24",X"6D",X"DD",X"EB",X"6D",X"55",X"55",
		X"49",X"49",X"2A",X"AD",X"DE",X"DD",X"DE",X"6E",X"B5",X"55",X"84",X"00",X"20",X"22",X"52",X"55",
		X"B5",X"56",X"6F",X"EB",X"F7",X"FF",X"FB",X"7B",X"B7",X"56",X"25",X"01",X"00",X"00",X"08",X"44",
		X"14",X"55",X"6B",X"DD",X"6D",X"DB",X"5A",X"B5",X"D6",X"5A",X"5B",X"AD",X"AA",X"A2",X"A4",X"52",
		X"A9",X"AA",X"6A",X"DB",X"7B",X"F7",X"76",X"AD",X"5A",X"95",X"24",X"49",X"8A",X"A4",X"54",X"B5",
		X"BD",X"B5",X"B5",X"6E",X"B7",X"7B",X"AB",X"55",X"20",X"10",X"04",X"01",X"02",X"21",X"24",X"4A",
		X"A9",X"52",X"52",X"24",X"92",X"CA",X"DA",X"F7",X"BF",X"FF",X"FF",X"FF",X"FB",X"BB",X"DB",X"AA",
		X"04",X"04",X"00",X"00",X"40",X"48",X"AA",X"AD",X"DD",X"DD",X"6E",X"5B",X"AB",X"4A",X"24",X"92",
		X"A4",X"D4",X"FE",X"FD",X"FF",X"BF",X"EF",X"6E",X"2D",X"89",X"40",X"00",X"82",X"10",X"89",X"52",
		X"B5",X"B6",X"5D",X"D7",X"AA",X"2A",X"4A",X"92",X"24",X"25",X"11",X"02",X"00",X"21",X"92",X"E2",
		X"FE",X"FF",X"FF",X"FF",X"EF",X"DE",X"AD",X"AA",X"14",X"22",X"00",X"00",X"40",X"10",X"A2",X"AA",
		X"BD",X"FF",X"FD",X"7D",X"BB",X"B5",X"52",X"10",X"00",X"10",X"84",X"94",X"AA",X"ED",X"EE",X"6E",
		X"EF",X"ED",X"6E",X"BB",X"5A",X"55",X"55",X"29",X"55",X"92",X"08",X"11",X"91",X"24",X"A9",X"76",
		X"FF",X"FB",X"BD",X"6D",X"2B",X"81",X"00",X"00",X"00",X"A1",X"A4",X"DA",X"EE",X"FB",X"7B",X"EF",
		X"AE",X"AB",X"55",X"95",X"A2",X"A4",X"4A",X"BB",X"D5",X"6A",X"2A",X"29",X"29",X"55",X"2A",X"53",
		X"49",X"12",X"02",X"10",X"89",X"54",X"A6",X"5A",X"AF",X"EF",X"F7",X"FE",X"7F",X"FF",X"DE",X"6D",
		X"53",X"25",X"01",X"01",X"00",X"00",X"41",X"24",X"D5",X"76",X"DF",X"FD",X"76",X"AB",X"55",X"A5",
		X"22",X"A5",X"AA",X"DE",X"DE",X"7D",X"77",X"6D",X"95",X"42",X"04",X"04",X"22",X"22",X"12",X"89",
		X"88",X"88",X"94",X"4A",X"BB",X"FF",X"FF",X"FF",X"BB",X"AD",X"4A",X"29",X"29",X"55",X"55",X"25",
		X"81",X"00",X"10",X"24",X"52",X"6A",X"DD",X"BD",X"EF",X"ED",X"76",X"B7",X"B5",X"6A",X"55",X"D5",
		X"B6",X"F7",X"DE",X"B6",X"5A",X"12",X"10",X"00",X"02",X"84",X"44",X"A9",X"5A",X"AB",X"DA",X"54",
		X"95",X"AA",X"DA",X"F6",X"FF",X"FF",X"EF",X"BB",X"AD",X"4A",X"02",X"01",X"80",X"40",X"10",X"22",
		X"92",X"A4",X"AA",X"6D",X"BF",X"FF",X"FE",X"7E",X"EF",X"B6",X"B5",X"AA",X"24",X"84",X"00",X"41",
		X"24",X"A9",X"6A",X"DB",X"7B",X"6F",X"6F",X"77",X"B7",X"6D",X"6B",X"55",X"85",X"00",X"00",X"00",
		X"00",X"88",X"28",X"D5",X"B6",X"77",X"EF",X"DD",X"AD",X"55",X"55",X"55",X"B5",X"B6",X"DD",X"76",
		X"6B",X"55",X"29",X"22",X"A1",X"54",X"55",X"DB",X"ED",X"DA",X"5A",X"55",X"84",X"20",X"80",X"00",
		X"02",X"11",X"49",X"55",X"B5",X"FD",X"FE",X"FF",X"FE",X"F7",X"DD",X"6D",X"55",X"55",X"42",X"44",
		X"08",X"11",X"49",X"6B",X"EF",X"F7",X"BD",X"6B",X"55",X"09",X"08",X"00",X"00",X"10",X"44",X"49",
		X"A9",X"D6",X"76",X"F7",X"FE",X"FD",X"EE",X"6E",X"5B",X"AB",X"54",X"22",X"89",X"88",X"A4",X"54",
		X"D5",X"5A",X"AF",X"BB",X"DD",X"BD",X"DD",X"AA",X"04",X"01",X"01",X"88",X"A4",X"5A",X"F7",X"76",
		X"5B",X"AB",X"2A",X"4A",X"89",X"24",X"91",X"94",X"94",X"4A",X"55",X"6D",X"D7",X"EB",X"DA",X"ED",
		X"FB",X"BE",X"77",X"D7",X"AA",X"84",X"40",X"10",X"22",X"A9",X"AA",X"76",X"77",X"7B",X"B5",X"2A",
		X"91",X"88",X"A4",X"54",X"ED",X"7B",X"EF",X"AE",X"AD",X"92",X"00",X"02",X"00",X"41",X"48",X"A4",
		X"AA",X"ED",X"F7",X"FB",X"7B",X"B7",X"AB",X"4A",X"22",X"91",X"94",X"AA",X"ED",X"BE",X"DF",X"FF",
		X"7D",X"6F",X"5B",X"55",X"12",X"08",X"00",X"01",X"00",X"00",X"42",X"48",X"5A",X"BB",X"DF",X"DF",
		X"F7",X"DD",X"B5",X"A6",X"4A",X"49",X"29",X"55",X"55",X"DB",X"BA",X"DD",X"B6",X"56",X"55",X"A1",
		X"88",X"08",X"21",X"04",X"04",X"81",X"20",X"44",X"94",X"AA",X"76",X"FF",X"F7",X"FF",X"DF",X"77",
		X"B7",X"B5",X"AA",X"2A",X"55",X"A9",X"AA",X"54",X"29",X"49",X"24",X"21",X"22",X"42",X"48",X"44",
		X"92",X"24",X"55",X"D5",X"DE",X"7B",X"EF",X"EE",X"D6",X"AA",X"92",X"10",X"11",X"91",X"24",X"55",
		X"D5",X"F6",X"EE",X"BB",X"77",X"77",X"6B",X"AD",X"AA",X"12",X"11",X"21",X"04",X"21",X"49",X"AA",
		X"6A",X"FB",X"EE",X"DD",X"ED",X"D6",X"B6",X"6A",X"55",X"AB",X"56",X"D5",X"AA",X"24",X"91",X"10",
		X"11",X"91",X"A4",X"6A",X"FB",X"F7",X"7B",X"77",X"6B",X"55",X"09",X"11",X"42",X"44",X"24",X"92",
		X"52",X"55",X"55",X"55",X"95",X"92",X"52",X"4A",X"A9",X"AA",X"AA",X"6A",X"DD",X"76",X"F7",X"BE",
		X"DF",X"BF",X"DF",X"BB",X"6D",X"55",X"55",X"42",X"84",X"10",X"91",X"A4",X"4A",X"55",X"55",X"55",
		X"B5",X"AA",X"AA",X"94",X"52",X"24",X"49",X"44",X"89",X"92",X"A2",X"A8",X"AA",X"FD",X"EE",X"DB",
		X"B6",X"5A",X"55",X"55",X"94",X"92",X"52",X"B5",X"BD",X"BB",X"DD",X"DA",X"AA",X"0A",X"89",X"A4",
		X"54",X"D5",X"7D",X"DF",X"77",X"77",X"B7",X"DD",X"B6",X"55",X"55",X"45",X"22",X"21",X"22",X"22",
		X"89",X"48",X"24",X"12",X"11",X"22",X"42",X"88",X"10",X"49",X"52",X"55",X"BB",X"DF",X"FF",X"FE",
		X"EF",X"FB",X"76",X"5B",X"55",X"95",X"24",X"12",X"49",X"49",X"A9",X"AA",X"B5",X"B6",X"AD",X"55",
		X"55",X"48",X"88",X"08",X"11",X"22",X"49",X"52",X"AA",X"AA",X"5A",X"6F",X"6B",X"6B",X"B5",X"AA",
		X"2A",X"55",X"AA",X"2A",X"55",X"55",X"AB",X"7D",X"DF",X"FB",X"EE",X"ED",X"B6",X"B5",X"AA",X"8A",
		X"48",X"49",X"A9",X"AA",X"AA",X"AA",X"AA",X"2A",X"09",X"21",X"88",X"48",X"A2",X"A4",X"54",X"AA",
		X"AA",X"EA",X"DE",X"F7",X"BD",X"77",X"BB",X"B6",X"AA",X"2A",X"12",X"25",X"49",X"24",X"A5",X"AA",
		X"EA",X"EE",X"EE",X"DE",X"6D",X"AF",X"56",X"95",X"20",X"04",X"21",X"22",X"95",X"6A",X"DB",X"DD",
		X"B6",X"DB",X"B6",X"6D",X"AB",X"2A",X"84",X"20",X"20",X"44",X"24",X"49",X"AA",X"6A",X"BD",X"77",
		X"EF",X"EE",X"B6",X"6D",X"D5",X"AA",X"AA",X"02",X"00",X"00",X"A0",X"7B",X"EF",X"EE",X"EA",X"FF",
		X"42",X"A2",X"B6",X"B6",X"70",X"11",X"82",X"80",X"80",X"28",X"35",X"BC",X"FF",X"FF",X"FF",X"87",
		X"00",X"09",X"89",X"44",X"25",X"01",X"00",X"00",X"4D",X"FD",X"F6",X"FF",X"FF",X"FF",X"FF",X"0B",
		X"00",X"00",X"C0",X"79",X"21",X"01",X"F4",X"FD",X"5B",X"A9",X"B3",X"00",X"FE",X"04",X"25",X"CC",
		X"DF",X"B6",X"56",X"49",X"90",X"54",X"F0",X"FF",X"FF",X"07",X"80",X"FD",X"03",X"13",X"C0",X"00",
		X"00",X"7E",X"01",X"28",X"BD",X"FF",X"FF",X"E3",X"FD",X"FF",X"5B",X"29",X"24",X"E0",X"17",X"40",
		X"FD",X"01",X"00",X"00",X"04",X"C2",X"7C",X"2B",X"49",X"70",X"ED",X"FF",X"FF",X"FF",X"FC",X"05",
		X"00",X"48",X"25",X"49",X"92",X"00",X"00",X"00",X"C0",X"BF",X"FF",X"FF",X"03",X"1C",X"FF",X"1F",
		X"1E",X"E2",X"1F",X"E9",X"57",X"00",X"00",X"38",X"9F",X"F7",X"FD",X"03",X"03",X"00",X"7C",X"FC",
		X"FF",X"45",X"00",X"FF",X"FF",X"0F",X"00",X"DA",X"03",X"FC",X"28",X"40",X"F5",X"EE",X"FF",X"FE",
		X"25",X"00",X"08",X"C7",X"41",X"7B",X"B7",X"AA",X"55",X"FD",X"17",X"0A",X"55",X"D2",X"67",X"00",
		X"10",X"29",X"18",X"FE",X"FF",X"EA",X"7D",X"9F",X"EA",X"7F",X"09",X"7C",X"3E",X"03",X"06",X"00",
		X"0A",X"40",X"00",X"80",X"FE",X"FF",X"FF",X"57",X"5A",X"F7",X"FF",X"FF",X"7F",X"8B",X"00",X"00",
		X"00",X"40",X"81",X"FF",X"A2",X"6B",X"FF",X"FD",X"01",X"00",X"FE",X"1F",X"00",X"D0",X"FF",X"FF",
		X"03",X"F0",X"41",X"FF",X"7F",X"55",X"04",X"00",X"E0",X"2A",X"44",X"ED",X"7F",X"2B",X"51",X"00",
		X"20",X"ED",X"FF",X"FF",X"DF",X"6F",X"6D",X"01",X"00",X"C0",X"F3",X"83",X"55",X"AD",X"84",X"3F",
		X"41",X"B6",X"FB",X"FD",X"03",X"60",X"04",X"80",X"A2",X"7F",X"FF",X"FF",X"87",X"10",X"0D",X"CE",
		X"F9",X"BF",X"16",X"08",X"00",X"00",X"90",X"FF",X"07",X"C0",X"FF",X"20",X"10",X"F5",X"FF",X"FF",
		X"44",X"D2",X"15",X"9E",X"FF",X"9F",X"23",X"05",X"00",X"40",X"3D",X"0E",X"1E",X"C0",X"1F",X"00",
		X"E8",X"F6",X"BF",X"BD",X"7C",X"70",X"66",X"10",X"3E",X"FF",X"FF",X"0A",X"05",X"E1",X"47",X"48",
		X"0F",X"41",X"0E",X"00",X"B0",X"07",X"A4",X"FD",X"FF",X"FF",X"FF",X"7F",X"DD",X"10",X"70",X"00",
		X"2F",X"E0",X"3F",X"01",X"40",X"A1",X"42",X"D5",X"56",X"00",X"00",X"7E",X"BD",X"7D",X"FB",X"BF",
		X"B3",X"FF",X"03",X"1E",X"87",X"00",X"00",X"4C",X"03",X"0B",X"F5",X"E0",X"75",X"B7",X"FD",X"DA",
		X"6B",X"1B",X"3F",X"4F",X"41",X"F0",X"04",X"00",X"00",X"C0",X"FB",X"4B",X"A4",X"EA",X"57",X"FF",
		X"F7",X"9F",X"59",X"C0",X"01",X"00",X"C0",X"03",X"70",X"C0",X"C3",X"5F",X"70",X"06",X"FA",X"FD",
		X"FD",X"E0",X"5C",X"CB",X"FF",X"FF",X"DF",X"AF",X"A0",X"00",X"02",X"00",X"12",X"00",X"80",X"FE",
		X"0F",X"45",X"F1",X"7F",X"7F",X"D1",X"FF",X"02",X"00",X"7F",X"FC",X"C1",X"BF",X"E0",X"8D",X"C7",
		X"FF",X"51",X"55",X"09",X"01",X"00",X"F0",X"7E",X"9B",X"A2",X"54",X"3F",X"7E",X"A9",X"3E",X"7F",
		X"FF",X"E1",X"03",X"FC",X"00",X"35",X"05",X"02",X"CC",X"1F",X"BF",X"EF",X"2F",X"00",X"00",X"AB",
		X"49",X"44",X"A2",X"3F",X"DE",X"FF",X"7F",X"D7",X"FF",X"08",X"80",X"80",X"5B",X"00",X"00",X"E8",
		X"7F",X"7F",X"97",X"00",X"C1",X"FF",X"FF",X"6A",X"05",X"00",X"00",X"B7",X"AF",X"F1",X"E7",X"7F",
		X"70",X"E0",X"C7",X"83",X"79",X"FC",X"7F",X"01",X"FC",X"D8",X"5A",X"05",X"00",X"00",X"42",X"ED",
		X"EF",X"F1",X"FF",X"F1",X"01",X"69",X"AD",X"B5",X"4A",X"EB",X"BE",X"D5",X"FF",X"28",X"24",X"25",
		X"29",X"02",X"18",X"04",X"50",X"D2",X"ED",X"FF",X"FB",X"FF",X"5F",X"FD",X"FB",X"1E",X"01",X"80",
		X"8A",X"00",X"00",X"40",X"F4",X"FF",X"FF",X"FF",X"95",X"24",X"ED",X"1F",X"EF",X"0F",X"25",X"41",
		X"00",X"00",X"10",X"08",X"E4",X"FF",X"FF",X"FF",X"FF",X"17",X"00",X"7F",X"70",X"00",X"E6",X"F7",
		X"FB",X"FF",X"7F",X"01",X"30",X"00",X"AC",X"5F",X"F5",X"A3",X"A4",X"F6",X"06",X"00",X"00",X"A4",
		X"FF",X"FF",X"FC",X"E3",X"F7",X"1B",X"70",X"01",X"00",X"F0",X"E7",X"FF",X"01",X"0D",X"14",X"80",
		X"AA",X"76",X"FD",X"FF",X"FF",X"7F",X"B5",X"01",X"00",X"00",X"E0",X"00",X"00",X"FC",X"3F",X"F8",
		X"FF",X"FF",X"C2",X"00",X"20",X"20",X"E2",X"AA",X"F8",X"FF",X"FF",X"2D",X"11",X"08",X"01",X"08",
		X"00",X"00",X"72",X"FB",X"FF",X"FF",X"7F",X"01",X"00",X"A0",X"80",X"4E",X"00",X"00",X"40",X"FE",
		X"3F",X"E0",X"20",X"68",X"3F",X"00",X"00",X"D4",X"54",X"F7",X"EB",X"EF",X"FF",X"0F",X"1C",X"00",
		X"00",X"01",X"00",X"00",X"FC",X"5F",X"CB",X"F6",X"FF",X"FF",X"8F",X"0F",X"00",X"00",X"14",X"00",
		X"EE",X"92",X"F6",X"FF",X"FF",X"4B",X"00",X"08",X"E4",X"03",X"00",X"50",X"6D",X"0E",X"FF",X"FF",
		X"4B",X"A8",X"FF",X"B7",X"55",X"34",X"00",X"00",X"00",X"D0",X"FF",X"7F",X"55",X"FB",X"FF",X"FF",
		X"FF",X"1B",X"00",X"FB",X"02",X"40",X"45",X"95",X"9F",X"E3",X"FF",X"FF",X"15",X"0A",X"55",X"15",
		X"19",X"A4",X"60",X"A0",X"B5",X"FF",X"FF",X"D7",X"FF",X"FF",X"FF",X"2E",X"02",X"00",X"00",X"00",
		X"00",X"EC",X"FA",X"FF",X"FF",X"3C",X"FF",X"FC",X"83",X"F3",X"F8",X"FC",X"C7",X"3E",X"5F",X"E4",
		X"17",X"00",X"00",X"D2",X"DB",X"2E",X"00",X"80",X"D7",X"FF",X"FF",X"FE",X"E1",X"A0",X"1F",X"7D",
		X"0D",X"00",X"F0",X"0F",X"FC",X"00",X"44",X"F2",X"00",X"02",X"E0",X"53",X"B5",X"F1",X"FF",X"FF",
		X"FF",X"01",X"80",X"BE",X"04",X"00",X"00",X"F8",X"7F",X"64",X"94",X"00",X"C7",X"FB",X"0F",X"04",
		X"10",X"1A",X"FC",X"BF",X"F4",X"FF",X"DF",X"55",X"20",X"70",X"00",X"06",X"A0",X"3F",X"02",X"8C",
		X"FE",X"C5",X"FF",X"FF",X"57",X"00",X"3D",X"08",X"02",X"15",X"00",X"00",X"80",X"FF",X"7B",X"FC",
		X"FE",X"FF",X"FF",X"0B",X"00",X"00",X"C0",X"FF",X"02",X"7F",X"C0",X"27",X"E0",X"0F",X"AC",X"7F",
		X"FC",X"02",X"06",X"FC",X"F1",X"DF",X"FF",X"6F",X"1D",X"0C",X"00",X"00",X"00",X"FA",X"FF",X"FF",
		X"43",X"75",X"01",X"70",X"7C",X"64",X"01",X"1A",X"04",X"EB",X"FF",X"87",X"FD",X"DF",X"08",X"1A",
		X"00",X"00",X"00",X"F8",X"FF",X"1C",X"FF",X"F7",X"FB",X"63",X"00",X"88",X"02",X"83",X"FF",X"FC",
		X"F7",X"80",X"0B",X"00",X"00",X"C1",X"C7",X"FF",X"FF",X"FF",X"50",X"84",X"BE",X"0A",X"A9",X"7D",
		X"41",X"34",X"56",X"4D",X"4B",X"04",X"02",X"50",X"F5",X"07",X"FD",X"F4",X"FF",X"FF",X"FF",X"05",
		X"00",X"00",X"A4",X"03",X"8B",X"EB",X"05",X"52",X"90",X"CF",X"EF",X"FF",X"FF",X"E8",X"1B",X"00",
		X"00",X"D0",X"FD",X"FF",X"01",X"71",X"01",X"00",X"EF",X"FF",X"BF",X"FA",X"0A",X"C0",X"FF",X"C0",
		X"8E",X"1E",X"00",X"FC",X"5E",X"11",X"10",X"E0",X"BA",X"3F",X"C0",X"1F",X"EA",X"E3",X"1F",X"E0",
		X"94",X"F0",X"FF",X"BF",X"0F",X"80",X"01",X"00",X"F8",X"FF",X"B3",X"DE",X"DA",X"00",X"00",X"00",
		X"41",X"F5",X"FD",X"FF",X"FF",X"7F",X"01",X"00",X"80",X"2C",X"FC",X"FF",X"5F",X"05",X"00",X"80",
		X"A8",X"55",X"FD",X"7F",X"FF",X"3F",X"07",X"70",X"00",X"00",X"20",X"F5",X"7E",X"F0",X"06",X"89",
		X"E8",X"FF",X"FC",X"5F",X"E0",X"F1",X"6F",X"50",X"85",X"4A",X"42",X"00",X"00",X"02",X"00",X"F5",
		X"FF",X"FF",X"7F",X"FF",X"3C",X"0C",X"00",X"00",X"04",X"28",X"7A",X"7D",X"BF",X"68",X"B1",X"43",
		X"92",X"E8",X"C1",X"00",X"00",X"00",X"F2",X"9F",X"FF",X"FF",X"FD",X"06",X"18",X"7E",X"2E",X"00",
		X"15",X"40",X"20",X"41",X"80",X"D4",X"FF",X"FF",X"3F",X"00",X"A0",X"EB",X"7F",X"3D",X"0B",X"F0",
		X"00",X"3B",X"FD",X"D1",X"A5",X"FF",X"D2",X"E1",X"1F",X"18",X"C0",X"01",X"00",X"88",X"8C",X"5F",
		X"FC",X"55",X"F5",X"EB",X"BB",X"2A",X"F0",X"7F",X"FE",X"7F",X"1C",X"00",X"00",X"01",X"02",X"80",
		X"00",X"A8",X"FE",X"FF",X"FF",X"9F",X"FF",X"78",X"09",X"10",X"80",X"E3",X"2F",X"02",X"FC",X"87",
		X"87",X"7B",X"00",X"00",X"01",X"8C",X"A7",X"51",X"37",X"A0",X"FF",X"3F",X"FF",X"FF",X"DF",X"05",
		X"A0",X"01",X"00",X"00",X"A0",X"C7",X"EF",X"E1",X"49",X"20",X"F0",X"FF",X"D6",X"FF",X"FF",X"DF",
		X"14",X"80",X"C3",X"00",X"00",X"A0",X"F4",X"7E",X"45",X"FE",X"1B",X"B0",X"B8",X"38",X"D0",X"7F",
		X"FF",X"3F",X"1D",X"00",X"40",X"7C",X"01",X"B4",X"EE",X"00",X"3B",X"AC",X"C2",X"01",X"FE",X"FF",
		X"FF",X"88",X"FF",X"FF",X"D5",X"01",X"E0",X"18",X"00",X"00",X"FA",X"3C",X"8E",X"03",X"3E",X"3E",
		X"FC",X"FF",X"BF",X"20",X"08",X"A0",X"FF",X"76",X"23",X"00",X"00",X"2B",X"3C",X"78",X"4E",X"40",
		X"17",X"18",X"40",X"D9",X"FF",X"DF",X"FF",X"56",X"8F",X"09",X"80",X"0F",X"74",X"7F",X"E6",X"C0",
		X"7F",X"00",X"00",X"0C",X"F8",X"FF",X"AF",X"E9",X"04",X"80",X"FA",X"AF",X"EA",X"FD",X"F7",X"AF",
		X"D7",X"05",X"00",X"00",X"00",X"21",X"FE",X"FF",X"CF",X"2A",X"01",X"F0",X"3C",X"FF",X"07",X"00",
		X"84",X"2D",X"DF",X"DA",X"3F",X"FC",X"5F",X"14",X"30",X"F0",X"7F",X"A8",X"7F",X"7E",X"38",X"C0",
		X"A5",X"86",X"08",X"3E",X"00",X"06",X"F8",X"FF",X"51",X"FA",X"FE",X"FB",X"DF",X"B7",X"40",X"00",
		X"00",X"F2",X"3E",X"9E",X"E9",X"03",X"80",X"FF",X"A1",X"7A",X"0D",X"84",X"15",X"E1",X"7F",X"37",
		X"5A",X"70",X"28",X"AE",X"FF",X"7F",X"BC",X"1F",X"4A",X"05",X"00",X"00",X"00",X"DA",X"E7",X"FB",
		X"3F",X"5C",X"94",X"F4",X"FF",X"0F",X"FD",X"F7",X"73",X"12",X"00",X"00",X"99",X"57",X"CF",X"07",
		X"2C",X"8E",X"01",X"00",X"FF",X"8E",X"D5",X"FF",X"FF",X"07",X"0E",X"00",X"FE",X"23",X"12",X"EB",
		X"FC",X"F9",X"A3",X"6C",X"A1",X"01",X"43",X"11",X"EA",X"FF",X"7F",X"F0",X"F0",X"80",X"90",X"03",
		X"BC",X"10",X"70",X"EF",X"FF",X"FF",X"42",X"4A",X"0F",X"C3",X"0A",X"6F",X"38",X"FC",X"E2",X"9F",
		X"4B",X"8A",X"C3",X"28",X"D5",X"0B",X"00",X"E0",X"27",X"8D",X"DE",X"EF",X"FF",X"FF",X"3F",X"01",
		X"00",X"00",X"BF",X"1F",X"1C",X"10",X"A4",X"2C",X"7F",X"FF",X"C9",X"A3",X"07",X"80",X"8F",X"F7",
		X"F9",X"F8",X"0D",X"C7",X"B5",X"FE",X"79",X"02",X"00",X"40",X"14",X"F8",X"1F",X"1E",X"7F",X"E0",
		X"81",X"1B",X"C2",X"EF",X"3F",X"01",X"61",X"71",X"E7",X"35",X"00",X"7C",X"96",X"FF",X"FC",X"0F",
		X"B4",X"FF",X"8B",X"00",X"40",X"CE",X"D7",X"0B",X"CB",X"0F",X"06",X"12",X"BA",X"54",X"0B",X"7D",
		X"FD",X"FF",X"FF",X"17",X"50",X"41",X"52",X"28",X"8E",X"41",X"30",X"0C",X"1E",X"8F",X"F8",X"EB",
		X"FF",X"7F",X"00",X"E0",X"01",X"FB",X"C1",X"07",X"DC",X"11",X"40",X"FD",X"FF",X"07",X"A1",X"7C",
		X"5E",X"EF",X"FF",X"02",X"10",X"C0",X"48",X"0D",X"F8",X"CA",X"FF",X"F7",X"B4",X"1D",X"01",X"00",
		X"C0",X"C7",X"F3",X"1F",X"BF",X"7E",X"17",X"F1",X"06",X"12",X"7C",X"E3",X"EF",X"3A",X"10",X"00",
		X"00",X"FD",X"F8",X"7B",X"D0",X"AF",X"0A",X"0A",X"98",X"DD",X"57",X"EB",X"FE",X"FF",X"AB",X"56",
		X"81",X"00",X"02",X"00",X"60",X"DD",X"FB",X"FF",X"1F",X"D5",X"7A",X"02",X"02",X"8E",X"8A",X"68",
		X"FD",X"FD",X"FE",X"BF",X"42",X"30",X"38",X"80",X"2D",X"96",X"F6",X"63",X"C0",X"FF",X"D2",X"5F",
		X"3F",X"2B",X"52",X"18",X"00",X"00",X"8C",X"C2",X"FE",X"FE",X"BE",X"CE",X"6F",X"01",X"98",X"C7",
		X"EB",X"25",X"1E",X"3E",X"43",X"49",X"05",X"B2",X"FC",X"F8",X"BF",X"D2",X"5A",X"4E",X"3F",X"01",
		X"00",X"AA",X"03",X"50",X"E3",X"F0",X"D7",X"FB",X"FD",X"FF",X"7F",X"5A",X"00",X"0A",X"20",X"00",
		X"F1",X"0E",X"3F",X"1F",X"A1",X"6E",X"04",X"30",X"FF",X"D5",X"FB",X"DF",X"2B",X"20",X"98",X"28",
		X"E0",X"EB",X"5D",X"97",X"76",X"D0",X"4A",X"04",X"06",X"84",X"E2",X"5B",X"FE",X"FF",X"FF",X"6B",
		X"07",X"10",X"03",X"04",X"C5",X"4E",X"F6",X"63",X"35",X"02",X"03",X"F8",X"07",X"A9",X"9F",X"FF",
		X"EA",X"FB",X"57",X"F4",X"02",X"00",X"30",X"DD",X"AA",X"F6",X"50",X"60",X"78",X"EC",X"97",X"07",
		X"F2",X"9F",X"FE",X"94",X"3E",X"F1",X"03",X"03",X"04",X"50",X"FD",X"E2",X"CF",X"1F",X"80",X"7A",
		X"C5",X"4F",X"3F",X"FC",X"03",X"0E",X"FC",X"60",X"5F",X"20",X"70",X"30",X"E0",X"F7",X"66",X"80",
		X"76",X"F7",X"07",X"4F",X"FD",X"FC",X"0F",X"42",X"D5",X"42",X"00",X"17",X"00",X"A4",X"FD",X"FF",
		X"E7",X"07",X"9F",X"12",X"00",X"57",X"35",X"77",X"D7",X"0F",X"3E",X"A9",X"AB",X"7A",X"50",X"60",
		X"01",X"38",X"F0",X"55",X"D7",X"F7",X"F5",X"DF",X"5F",X"45",X"80",X"05",X"C0",X"7E",X"01",X"8B",
		X"F4",X"D0",X"56",X"3F",X"20",X"A5",X"00",X"F4",X"DF",X"7F",X"E3",X"57",X"0A",X"5F",X"FA",X"AB",
		X"07",X"54",X"49",X"10",X"00",X"20",X"D0",X"FB",X"FF",X"FB",X"0D",X"0E",X"78",X"F8",X"AF",X"A4",
		X"50",X"A9",X"FE",X"C0",X"32",X"4C",X"15",X"50",X"F4",X"FF",X"9F",X"B5",X"60",X"04",X"44",X"EE",
		X"8E",X"BE",X"FC",X"A8",X"00",X"F8",X"C0",X"7E",X"EC",X"BF",X"C2",X"40",X"D5",X"FD",X"F8",X"B0",
		X"0E",X"04",X"48",X"C6",X"87",X"FB",X"2F",X"1C",X"38",X"EF",X"3F",X"0C",X"D1",X"C3",X"F9",X"3F",
		X"80",X"0E",X"B1",X"46",X"80",X"87",X"67",X"F9",X"F1",X"AF",X"20",X"74",X"75",X"BD",X"E0",X"43",
		X"B7",X"4A",X"21",X"38",X"80",X"69",X"FF",X"5F",X"FE",X"08",X"02",X"3C",X"3E",X"8B",X"6A",X"7D",
		X"70",X"E0",X"11",X"FB",X"F7",X"36",X"E0",X"D5",X"72",X"FA",X"36",X"55",X"00",X"00",X"80",X"EB",
		X"7F",X"5B",X"60",X"D1",X"5E",X"FD",X"3F",X"C1",X"22",X"C2",X"D5",X"5F",X"2F",X"DA",X"57",X"0B",
		X"12",X"00",X"67",X"40",X"1F",X"FC",X"2C",X"66",X"C9",X"67",X"FF",X"09",X"38",X"16",X"65",X"E3",
		X"7F",X"ED",X"F0",X"A9",X"C0",X"A0",X"A3",X"5D",X"57",X"08",X"C7",X"06",X"49",X"60",X"68",X"A3",
		X"FA",X"FF",X"AF",X"FF",X"55",X"80",X"95",X"D0",X"07",X"2C",X"59",X"00",X"F2",X"C0",X"FB",X"4A",
		X"7F",X"DE",X"FB",X"A9",X"0A",X"E0",X"00",X"C2",X"27",X"7F",X"6A",X"2B",X"7E",X"8C",X"B7",X"0B",
		X"00",X"7E",X"F0",X"45",X"FB",X"2F",X"51",X"54",X"F8",X"D7",X"05",X"00",X"A2",X"F1",X"E1",X"BD",
		X"A0",X"B6",X"7A",X"FD",X"77",X"2F",X"52",X"C0",X"40",X"E8",X"DF",X"CB",X"80",X"B0",X"F6",X"AF",
		X"11",X"10",X"FA",X"03",X"7C",X"62",X"53",X"7E",X"BC",X"6B",X"87",X"02",X"F8",X"D0",X"FE",X"D7",
		X"00",X"8F",X"5F",X"B5",X"05",X"80",X"D2",X"47",X"E9",X"03",X"A1",X"92",X"9F",X"E3",X"BF",X"C2",
		X"29",X"B0",X"7E",X"B1",X"FF",X"82",X"C1",X"39",X"EC",X"F4",X"C0",X"4F",X"00",X"CE",X"80",X"F3",
		X"3E",X"F6",X"E3",X"22",X"FC",X"F8",X"1E",X"AE",X"FA",X"55",X"12",X"08",X"C0",X"83",X"16",X"47",
		X"FF",X"2B",X"A8",X"83",X"F6",X"5F",X"50",X"12",X"AF",X"22",X"E2",X"BF",X"45",X"56",X"C5",X"87",
		X"7E",X"50",X"10",X"BC",X"C4",X"3F",X"AE",X"5D",X"4C",X"30",X"1D",X"C1",X"E1",X"E7",X"05",X"7E",
		X"60",X"15",X"FA",X"F0",X"FA",X"F1",X"58",X"24",X"85",X"FF",X"F3",X"1D",X"30",X"1E",X"04",X"92",
		X"8A",X"9E",X"00",X"2A",X"BA",X"BE",X"FA",X"81",X"5F",X"DF",X"74",X"7F",X"5F",X"BA",X"80",X"02",
		X"41",X"ED",X"44",X"2B",X"4F",X"A0",X"A4",X"5F",X"BD",X"C9",X"BF",X"05",X"80",X"83",X"56",X"FB",
		X"89",X"C2",X"BF",X"AE",X"49",X"BF",X"2E",X"00",X"A5",X"92",X"54",X"11",X"16",X"F7",X"FF",X"DD",
		X"F0",X"80",X"83",X"9E",X"63",X"30",X"D0",X"75",X"FF",X"F1",X"2A",X"11",X"14",X"FD",X"A8",X"BF",
		X"5A",X"05",X"08",X"54",X"AB",X"BF",X"1E",X"A1",X"40",X"1E",X"20",X"F5",X"B7",X"57",X"6D",X"D5",
		X"8B",X"FA",X"0D",X"D0",X"07",X"59",X"D1",X"1A",X"DD",X"96",X"E8",X"0B",X"97",X"5F",X"09",X"08",
		X"21",X"DC",X"96",X"1C",X"B4",X"9A",X"BD",X"FE",X"FF",X"1F",X"BE",X"10",X"04",X"95",X"D0",X"F5",
		X"83",X"0B",X"10",X"1E",X"D3",X"6A",X"25",X"B2",X"FD",X"F3",X"21",X"37",X"BF",X"54",X"40",X"16",
		X"3C",X"52",X"2E",X"83",X"74",X"D2",X"9B",X"BB",X"AA",X"7E",X"BF",X"8E",X"41",X"01",X"1B",X"A3",
		X"64",X"B9",X"AE",X"E0",X"87",X"BF",X"1A",X"A1",X"C7",X"3F",X"6C",X"B5",X"0F",X"1C",X"8F",X"89",
		X"23",X"50",X"43",X"00",X"3C",X"55",X"70",X"2B",X"7C",X"FD",X"CF",X"3F",X"C2",X"D6",X"0A",X"7D",
		X"90",X"02",X"5D",X"AD",X"F0",X"45",X"83",X"6A",X"45",X"55",X"8A",X"B5",X"B3",X"3E",X"FD",X"F7",
		X"9F",X"0B",X"70",X"45",X"02",X"50",X"D5",X"AB",X"6A",X"7B",X"52",X"52",X"7F",X"E1",X"2F",X"15",
		X"A6",X"01",X"02",X"AF",X"62",X"01",X"5F",X"B7",X"EA",X"AA",X"7E",X"65",X"55",X"10",X"E8",X"F8",
		X"F8",X"06",X"C7",X"2F",X"87",X"42",X"FB",X"A9",X"0B",X"70",X"40",X"DB",X"57",X"7B",X"41",X"0F",
		X"97",X"2B",X"F2",X"A3",X"31",X"E0",X"6D",X"70",X"D0",X"D5",X"45",X"53",X"A5",X"FB",X"7E",X"6E",
		X"29",X"A8",X"00",X"CE",X"41",X"B7",X"5A",X"BD",X"00",X"55",X"6F",X"A0",X"5A",X"7D",X"E1",X"AF",
		X"0F",X"AA",X"85",X"87",X"4F",X"32",X"2C",X"0B",X"EA",X"A2",X"42",X"2B",X"62",X"AF",X"0F",X"5F",
		X"A1",X"D9",X"BE",X"5C",X"B5",X"0B",X"2F",X"D2",X"8F",X"2D",X"E4",X"E1",X"80",X"41",X"69",X"B1",
		X"8A",X"8A",X"DA",X"C3",X"7F",X"DA",X"56",X"D7",X"55",X"D8",X"A1",X"04",X"2A",X"D0",X"4A",X"95",
		X"DE",X"EB",X"8D",X"DB",X"A5",X"10",X"15",X"12",X"54",X"5D",X"FC",X"7C",X"75",X"4D",X"AF",X"B4",
		X"2C",X"3A",X"B0",X"D1",X"26",X"16",X"FA",X"C0",X"2F",X"FD",X"C0",X"0B",X"A4",X"6B",X"10",X"7A",
		X"81",X"7E",X"D0",X"B9",X"8E",X"6F",X"E9",X"BB",X"A2",X"DE",X"02",X"4A",X"59",X"55",X"84",X"AE",
		X"58",X"55",X"4B",X"5E",X"21",X"2A",X"5D",X"5E",X"AB",X"5F",X"B5",X"C0",X"E8",X"51",X"7A",X"61",
		X"3F",X"1A",X"C6",X"A8",X"7E",X"10",X"85",X"87",X"47",X"1E",X"3F",X"2E",X"1F",X"F8",X"70",X"8B",
		X"7D",X"8D",X"F0",X"19",X"17",X"0F",X"E8",X"50",X"45",X"29",X"A5",X"A8",X"EB",X"D9",X"D3",X"94",
		X"AD",X"FE",X"3F",X"3C",X"D4",X"29",X"50",X"54",X"49",X"B9",X"C0",X"51",X"C1",X"33",X"DE",X"72",
		X"EF",X"15",X"E3",X"DA",X"44",X"57",X"48",X"0E",X"71",X"DC",X"75",X"59",X"5F",X"A8",X"41",X"3D",
		X"14",X"95",X"A2",X"A9",X"74",X"BA",X"6F",X"FD",X"BA",X"A8",X"0B",X"54",X"A8",X"50",X"0F",X"3E",
		X"B4",X"4A",X"56",X"D0",X"D2",X"5A",X"5F",X"E9",X"AA",X"AE",X"F2",X"C1",X"82",X"64",X"AD",X"86",
		X"1E",X"54",X"7F",X"1D",X"97",X"AA",X"17",X"5E",X"38",X"02",X"27",X"09",X"6A",X"75",X"5F",X"19",
		X"EE",X"4B",X"94",X"EB",X"B2",X"AA",X"76",X"6B",X"89",X"83",X"42",X"D1",X"83",X"AB",X"52",X"A9",
		X"17",X"AF",X"4A",X"08",X"9A",X"AA",X"F6",X"5E",X"7D",X"95",X"AA",X"E2",X"F0",X"AD",X"88",X"2A",
		X"74",X"A5",X"1E",X"94",X"AA",X"92",X"AA",X"F4",X"EB",X"67",X"79",X"E0",X"C2",X"06",X"8F",X"E3",
		X"12",X"95",X"B5",X"1B",X"96",X"BA",X"48",X"25",X"55",X"AD",X"F4",X"AB",X"06",X"DE",X"A2",X"28",
		X"75",X"77",X"A5",X"2D",X"70",X"D1",X"2B",X"EF",X"52",X"81",X"1E",X"74",X"A5",X"0B",X"0F",X"56",
		X"45",X"55",X"9D",X"9E",X"56",X"AB",X"4A",X"A1",X"8A",X"74",X"F9",X"55",X"4F",X"16",X"54",X"45",
		X"BF",X"5A",X"A2",X"A4",X"76",X"74",X"AA",X"0A",X"54",X"D1",X"A5",X"8D",X"F6",X"A5",X"4B",X"5D",
		X"E4",X"55",X"9D",X"92",X"CD",X"0B",X"B4",X"14",X"CA",X"30",X"B5",X"F4",X"24",X"AD",X"EC",X"F2",
		X"AF",X"6C",X"0D",X"A5",X"2A",X"48",X"AB",X"52",X"D5",X"79",X"95",X"5E",X"55",X"D1",X"11",X"16",
		X"6D",X"95",X"96",X"F5",X"F2",X"C1",X"2B",X"EA",X"52",X"24",X"F5",X"50",X"A9",X"1E",X"7A",X"61",
		X"B7",X"0A",X"B6",X"52",X"55",X"D5",X"D5",X"85",X"B7",X"A5",X"C0",X"85",X"4D",X"55",X"95",X"2D",
		X"3D",X"7A",X"55",X"AB",X"38",X"AA",X"4A",X"55",X"EA",X"94",X"42",X"56",X"B1",X"EA",X"A8",X"F5",
		X"D5",X"A6",X"5A",X"52",X"2F",X"0E",X"12",X"A1",X"6A",X"5B",X"D4",X"A2",X"A7",X"6F",X"17",X"AB",
		X"2A",X"D8",X"51",X"55",X"75",X"C8",X"8A",X"F5",X"D5",X"85",X"2A",X"2D",X"A9",X"82",X"AB",X"5A",
		X"D5",X"95",X"DF",X"52",X"31",X"54",X"2D",X"B1",X"89",X"AB",X"F4",X"8A",X"AB",X"5E",X"22",X"45",
		X"AB",X"6A",X"D1",X"AA",X"83",X"CB",X"C3",X"47",X"E1",X"41",X"87",X"A3",X"C3",X"47",X"97",X"A5",
		X"57",X"D2",X"75",X"55",X"C5",X"9A",X"4A",X"51",X"A5",X"52",X"B4",X"72",X"5B",X"55",X"5D",X"54",
		X"97",X"52",X"72",X"89",X"7B",X"AB",X"B5",X"AA",X"57",X"55",X"D0",X"C8",X"41",X"55",X"15",X"47",
		X"8B",X"AA",X"95",X"5A",X"1D",X"A1",X"55",X"2D",X"E5",X"A9",X"FE",X"0A",X"A3",X"57",X"54",X"D1",
		X"1D",X"1E",X"C7",X"43",X"55",X"AC",X"AA",X"A3",X"4B",X"55",X"D5",X"45",X"8D",X"5A",X"55",X"5D",
		X"A5",X"B4",X"AA",X"2A",X"55",X"55",X"A5",X"2A",X"2A",X"51",X"15",X"6D",X"A9",X"FA",X"A0",X"8A",
		X"5A",X"D5",X"5D",X"D7",X"E3",X"54",X"AD",X"56",X"AB",X"3A",X"34",X"A5",X"45",X"2D",X"51",X"A1",
		X"4A",X"4A",X"D3",X"95",X"5D",X"5E",X"A5",X"BD",X"5A",X"DB",X"44",X"55",X"55",X"55",X"A2",X"D4",
		X"29",X"51",X"91",X"46",X"AA",X"4A",X"54",X"DD",X"E9",X"DB",X"3A",X"DB",X"5A",X"55",X"45",X"52",
		X"29",X"AE",X"B4",X"AA",X"8F",X"A8",X"C8",X"4C",X"97",X"D0",X"65",X"55",X"59",X"7D",X"D5",X"AB",
		X"55",X"55",X"A8",X"6A",X"55",X"29",X"85",X"2A",X"55",X"A5",X"2A",X"AE",X"D4",X"CA",X"AF",X"B6",
		X"D5",X"55",X"51",X"68",X"94",X"0E",X"AD",X"EA",X"55",X"0B",X"AD",X"52",X"95",X"5E",X"D5",X"52",
		X"95",X"AA",X"A4",X"E3",X"2A",X"55",X"55",X"8F",X"AA",X"A8",X"48",X"AD",X"3E",X"7A",X"AD",X"2A",
		X"BD",X"E8",X"4A",X"25",X"A5",X"AA",X"2A",X"D4",X"52",X"A3",X"16",X"CA",X"C3",X"87",X"1F",X"1E",
		X"BE",X"44",X"1F",X"87",X"E3",X"71",X"E8",X"F0",X"B0",X"16",X"4D",X"1D",X"0F",X"75",X"B9",X"94",
		X"CA",X"A6",X"97",X"16",X"6A",X"75",X"A1",X"55",X"55",X"92",X"56",X"AB",X"54",X"75",X"19",X"7A",
		X"D4",X"15",X"5E",X"74",X"55",X"1C",X"BD",X"F8",X"D0",X"89",X"A5",X"D2",X"52",X"B5",X"54",X"7A",
		X"1C",X"A5",X"5A",X"1D",X"D5",X"75",X"55",X"34",X"BD",X"54",X"45",X"4B",X"A5",X"6A",X"79",X"71",
		X"D4",X"51",X"AB",X"4A",X"55",X"A5",X"E2",X"AA",X"4A",X"AB",X"A6",X"4A",X"5F",X"AB",X"4A",X"45",
		X"8F",X"16",X"55",X"69",X"69",X"55",X"AD",X"52",X"2D",X"54",X"85",X"A3",X"D6",X"A2",X"55",X"D5",
		X"74",X"F4",X"6A",X"AB",X"52",X"95",X"8A",X"AA",X"56",X"C3",X"AF",X"4A",X"AA",X"AA",X"54",X"59",
		X"A1",X"72",X"55",X"D5",X"2E",X"1D",X"5D",X"92",X"92",X"36",X"BD",X"52",X"6F",X"75",X"45",X"45",
		X"55",X"AA",X"A4",X"DA",X"D2",X"D2",X"D2",X"96",X"74",X"55",X"16",X"2A",X"51",X"85",X"1D",X"7D",
		X"57",X"AD",X"AA",X"95",X"AA",X"5B",X"A8",X"5A",X"45",X"95",X"54",X"D2",X"85",X"56",X"4F",X"57",
		X"55",X"F4",X"E1",X"45",X"B5",X"16",X"27",X"4B",X"9D",X"AA",X"A5",X"AA",X"54",X"A5",X"96",X"56",
		X"55",X"A5",X"76",X"4A",X"2A",X"55",X"35",X"AC",X"AA",X"AA",X"B5",X"D2",X"6F",X"2D",X"5D",X"54",
		X"54",X"AA",X"6A",X"55",X"45",X"6B",X"A8",X"51",X"55",X"5F",X"74",X"AB",X"5A",X"A8",X"51",X"55",
		X"4D",X"D4",X"D2",X"55",X"6A",X"77",X"AB",X"EA",X"56",X"A4",X"0A",X"AC",X"AA",X"42",X"95",X"56",
		X"B5",X"D5",X"5B",X"55",X"22",X"AD",X"54",X"F5",X"2B",X"5B",X"54",X"15",X"8D",X"BA",X"EA",X"16",
		X"A5",X"AA",X"D2",X"A5",X"56",X"A9",X"4A",X"A5",X"AA",X"F2",X"95",X"5E",X"9A",X"A2",X"52",X"A5",
		X"55",X"A7",X"5A",X"A8",X"D4",X"4A",X"AD",X"5A",X"5A",X"9D",X"AA",X"4B",X"95",X"AA",X"A8",X"A8",
		X"2A",X"7D",X"AA",X"54",X"AD",X"2A",X"41",X"A5",X"AA",X"6A",X"AB",X"2E",X"55",X"55",X"65",X"55",
		X"D4",X"AA",X"95",X"A4",X"AA",X"55",X"5D",X"68",X"51",X"69",X"55",X"5D",X"5D",X"5D",X"51",X"55",
		X"55",X"55",X"D5",X"4A",X"2D",X"6A",X"A9",X"AA",X"54",X"AB",X"AB",X"1E",X"55",X"2F",X"4A",X"BA",
		X"54",X"55",X"55",X"55",X"53",X"AD",X"B2",X"B4",X"50",X"2D",X"D5",X"16",X"55",X"55",X"55",X"D5",
		X"55",X"55",X"D5",X"FA",X"2A",X"55",X"68",X"A9",X"96",X"D2",X"52",X"55",X"55",X"D5",X"55",X"55",
		X"55",X"15",X"95",X"D6",X"6A",X"A9",X"96",X"54",X"55",X"AD",X"AB",X"AA",X"50",X"A1",X"56",X"55",
		X"AB",X"AA",X"AA",X"6A",X"55",X"2B",X"15",X"69",X"D5",X"52",X"A9",X"2A",X"55",X"BD",X"6A",X"55",
		X"55",X"55",X"AA",X"52",X"55",X"55",X"A9",X"56",X"D5",X"AA",X"AB",X"2F",X"55",X"D4",X"A2",X"52",
		X"A9",X"AA",X"AA",X"2E",X"55",X"55",X"69",X"55",X"D5",X"55",X"55",X"D4",X"AA",X"55",X"95",X"AA",
		X"12",X"55",X"69",X"D5",X"AB",X"AA",X"A8",X"52",X"55",X"BA",X"AA",X"15",X"55",X"B5",X"AB",X"4A",
		X"55",X"54",X"5D",X"5A",X"B5",X"44",X"95",X"AE",X"AA",X"4A",X"B5",X"AA",X"52",X"25",X"B5",X"AA",
		X"AA",X"AE",X"6A",X"D5",X"4B",X"55",X"A8",X"AA",X"16",X"55",X"55",X"95",X"DA",X"EA",X"2B",X"55",
		X"95",X"AA",X"A2",X"16",X"5D",X"A5",X"55",X"55",X"7F",X"FC",X"FF",X"FF",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"C0",X"60",X"30",X"20",X"00",
		X"04",X"00",X"00",X"F8",X"F3",X"FC",X"FF",X"FB",X"0F",X"00",X"00",X"CF",X"FF",X"FF",X"00",X"30",
		X"70",X"E8",X"FF",X"01",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"01",X"00",
		X"A0",X"E1",X"7F",X"FE",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"FE",X"01",X"F0",X"5F",X"D5",
		X"81",X"03",X"FE",X"00",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"22",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"2F",X"FC",X"FF",X"FF",X"FF",X"03",X"00",X"7C",X"02",X"00",X"E0",
		X"FF",X"FF",X"C3",X"00",X"1E",X"00",X"00",X"00",X"F4",X"FF",X"FD",X"BF",X"FF",X"FF",X"0F",X"84",
		X"C0",X"00",X"00",X"00",X"CE",X"F9",X"FF",X"FF",X"00",X"00",X"00",X"72",X"E0",X"FF",X"FF",X"FF",
		X"01",X"00",X"00",X"80",X"FF",X"0F",X"70",X"00",X"00",X"C0",X"FF",X"FF",X"FF",X"07",X"C0",X"01",
		X"00",X"00",X"BD",X"FF",X"C7",X"EF",X"7F",X"00",X"F8",X"7F",X"05",X"00",X"38",X"00",X"00",X"00",
		X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"FC",X"5F",X"C1",X"01",X"00",X"00",X"00",X"00",X"C0",X"FF",
		X"FF",X"FF",X"02",X"00",X"F0",X"FF",X"7F",X"01",X"00",X"28",X"00",X"00",X"00",X"E0",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"2F",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"80",X"07",X"00",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"C3",X"0F",X"80",X"00",X"07",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E8",X"1F",X"86",X"87",X"E7",X"3F",X"7F",X"60",X"EE",X"FF",X"FF",X"FF",X"FF",X"07",X"40",
		X"00",X"20",X"30",X"60",X"F0",X"07",X"00",X"00",X"00",X"00",X"02",X"00",X"82",X"E3",X"FD",X"3F",
		X"8E",X"FF",X"FF",X"FF",X"FF",X"07",X"00",X"FF",X"FF",X"FF",X"0F",X"00",X"00",X"00",X"80",X"FF",
		X"07",X"00",X"78",X"00",X"00",X"00",X"00",X"41",X"1F",X"7F",X"3C",X"FF",X"FF",X"FF",X"19",X"F0",
		X"E1",X"C0",X"F9",X"77",X"FE",X"FF",X"3E",X"8F",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"04",
		X"07",X"CF",X"EF",X"3F",X"80",X"C7",X"CF",X"CF",X"63",X"70",X"03",X"FF",X"F3",X"E3",X"FF",X"FF",
		X"F3",X"01",X"06",X"00",X"83",X"E7",X"01",X"00",X"F8",X"FF",X"1F",X"C3",X"00",X"60",X"C0",X"F0",
		X"CD",X"F3",X"EF",X"0F",X"CE",X"FF",X"FF",X"FF",X"00",X"00",X"30",X"40",X"FD",X"05",X"FF",X"FF",
		X"FF",X"3F",X"00",X"00",X"00",X"80",X"FE",X"FB",X"FF",X"1F",X"7F",X"00",X"FF",X"CF",X"0F",X"18",
		X"0C",X"03",X"F0",X"83",X"EF",X"C7",X"CF",X"E3",X"FF",X"FF",X"FD",X"7F",X"00",X"38",X"E2",X"E0",
		X"80",X"01",X"06",X"C0",X"FF",X"1F",X"00",X"00",X"00",X"F8",X"FF",X"F1",X"EF",X"BF",X"FF",X"0D",
		X"00",X"00",X"00",X"F8",X"F3",X"E7",X"FF",X"FF",X"02",X"00",X"00",X"00",X"FE",X"FF",X"07",X"FF",
		X"FF",X"7F",X"C7",X"00",X"07",X"00",X"00",X"80",X"87",X"7F",X"BE",X"FF",X"FF",X"1F",X"0C",X"0C",
		X"80",X"40",X"F8",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F8",X"E3",X"DF",X"FB",X"BF",X"1B",X"00",
		X"10",X"16",X"4E",X"0E",X"43",X"38",X"FC",X"38",X"78",X"9C",X"FF",X"FF",X"7F",X"1E",X"00",X"00",
		X"00",X"FE",X"FF",X"FF",X"1F",X"F3",X"07",X"00",X"C0",X"FF",X"9F",X"80",X"0F",X"00",X"00",X"00",
		X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"83",X"FF",X"FF",X"07",X"00",X"00",X"06",X"00",X"00",X"00",
		X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"8B",X"01",X"86",X"6A",X"3F",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"0F",X"03",X"8C",X"FF",X"7F",X"63",X"29",X"A9",X"2A",X"45",X"40",X"70",X"1E",X"09",
		X"00",X"00",X"00",X"08",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"27",X"0E",X"00",X"60",X"FF",X"FF",
		X"FF",X"FF",X"8F",X"FF",X"7F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"BF",X"FF",
		X"FF",X"FF",X"CB",X"FF",X"FF",X"DF",X"09",X"00",X"C0",X"30",X"84",X"7F",X"E0",X"DD",X"E7",X"0F",
		X"0E",X"C7",X"CF",X"C7",X"00",X"00",X"00",X"70",X"C1",X"CF",X"F1",X"1C",X"1E",X"1C",X"00",X"CF",
		X"39",X"07",X"07",X"1F",X"77",X"3C",X"3F",X"B8",X"71",X"B0",X"0F",X"E0",X"EF",X"FF",X"F1",X"03",
		X"0F",X"E0",X"00",X"00",X"00",X"F0",X"7C",X"FF",X"78",X"C0",X"81",X"FF",X"FF",X"1F",X"80",X"01",
		X"00",X"04",X"FF",X"FF",X"FF",X"FB",X"FF",X"FF",X"3D",X"80",X"07",X"00",X"00",X"00",X"00",X"B0",
		X"E3",X"C7",X"F3",X"FF",X"FF",X"F0",X"80",X"01",X"01",X"8C",X"FF",X"FE",X"FC",X"3B",X"3E",X"7C",
		X"78",X"1C",X"08",X"00",X"82",X"8F",X"1F",X"F7",X"61",X"00",X"99",X"FF",X"C6",X"83",X"19",X"FC",
		X"00",X"3E",X"F9",X"C0",X"87",X"00",X"00",X"E0",X"7F",X"FE",X"F8",X"3F",X"00",X"00",X"00",X"C0",
		X"FF",X"FB",X"8F",X"FF",X"FF",X"3F",X"38",X"0C",X"37",X"7C",X"0E",X"00",X"00",X"00",X"00",X"FF",
		X"F7",X"C7",X"CF",X"FB",X"CF",X"0D",X"02",X"03",X"02",X"00",X"60",X"F0",X"77",X"CF",X"07",X"0C",
		X"10",X"E7",X"3F",X"38",X"FE",X"3F",X"1E",X"0E",X"1C",X"F1",X"03",X"7F",X"38",X"87",X"DF",X"F1",
		X"C7",X"31",X"08",X"70",X"C0",X"E3",X"C8",X"9F",X"07",X"07",X"00",X"80",X"83",X"FF",X"0B",X"E3",
		X"39",X"FF",X"3F",X"C3",X"31",X"84",X"21",X"98",X"C3",X"70",X"02",X"FE",X"F0",X"FF",X"FF",X"3E",
		X"01",X"80",X"00",X"EE",X"FE",X"F1",X"3F",X"E0",X"BF",X"FF",X"7F",X"1F",X"00",X"00",X"00",X"00",
		X"F4",X"E0",X"FF",X"FF",X"FF",X"67",X"08",X"38",X"70",X"00",X"00",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"10",X"C0",X"01",X"00",X"00",X"20",X"58",X"55",X"2A",X"F0",X"E7",X"FF",X"31",X"64",X"38",
		X"38",X"CC",X"FF",X"3F",X"3F",X"04",X"00",X"E0",X"FF",X"FF",X"FF",X"1F",X"04",X"00",X"00",X"00",
		X"00",X"34",X"7E",X"FE",X"8F",X"07",X"C7",X"FD",X"FF",X"BF",X"00",X"00",X"00",X"E0",X"FF",X"F7",
		X"FF",X"FF",X"1F",X"E0",X"FF",X"02",X"00",X"06",X"00",X"00",X"00",X"00",X"88",X"FF",X"FF",X"38",
		X"E7",X"FF",X"3F",X"0F",X"00",X"00",X"E8",X"FE",X"82",X"D4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"C3",X"01",X"C4",X"03",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"7F",X"FF",X"01",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"2B",X"00",X"7C",X"03",X"00",X"00",X"18",X"00",X"00",
		X"00",X"82",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7B",X"18",X"F0",X"7F",X"1E",X"00",X"00",
		X"00",X"00",X"00",X"EF",X"FF",X"47",X"70",X"00",X"00",X"90",X"7F",X"FF",X"FF",X"FF",X"3F",X"9E",
		X"1F",X"00",X"00",X"00",X"80",X"FF",X"56",X"E9",X"19",X"30",X"C0",X"FF",X"0F",X"06",X"FE",X"FB",
		X"3F",X"FC",X"FF",X"FF",X"FF",X"07",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"07",
		X"F8",X"FF",X"BF",X"00",X"00",X"00",X"00",X"E0",X"07",X"04",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"44",X"1C",X"7F",X"CF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"03",X"00",X"01",X"08",X"00",X"03",X"08",X"00",X"08",X"19",
		X"70",X"FE",X"FF",X"7B",X"3E",X"C0",X"C1",X"FF",X"FF",X"FF",X"07",X"00",X"00",X"D0",X"FF",X"FF",
		X"7F",X"E0",X"FF",X"BF",X"70",X"00",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FF",X"BF",X"EF",X"FF",
		X"FF",X"7F",X"00",X"00",X"00",X"F8",X"E7",X"FF",X"30",X"F0",X"39",X"0C",X"EC",X"38",X"FF",X"FF",
		X"BB",X"00",X"10",X"38",X"18",X"04",X"E0",X"E0",X"60",X"DC",X"EF",X"01",X"3B",X"9E",X"FF",X"FE",
		X"FF",X"07",X"00",X"00",X"E8",X"0F",X"FF",X"F8",X"3F",X"1E",X"87",X"01",X"3C",X"04",X"00",X"00",
		X"60",X"03",X"07",X"E7",X"FD",X"FF",X"03",X"C6",X"E1",X"1F",X"00",X"FE",X"FF",X"FF",X"FF",X"0F",
		X"10",X"00",X"78",X"07",X"B0",X"FF",X"FF",X"FF",X"8F",X"C3",X"FF",X"FF",X"03",X"00",X"00",X"00",
		X"00",X"18",X"EE",X"73",X"7C",X"FF",X"FF",X"39",X"04",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"3F",X"00",X"00",X"00",X"C0",X"3F",X"FE",X"F7",X"FF",X"0F",X"00",X"C0",X"BF",X"09",X"00",X"00",
		X"C0",X"03",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"7F",X"0E",X"00",X"FF",X"01",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"FE",X"BF",X"20",X"44",
		X"10",X"00",X"FF",X"03",X"00",X"18",X"04",X"06",X"C3",X"40",X"FC",X"7F",X"3C",X"FC",X"FF",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"07",X"00",X"A8",X"ED",X"B6",X"24",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"19",X"FC",X"FF",X"E7",X"79",X"3C",X"38",X"FC",X"FF",X"FF",X"FF",X"7F",X"FF",
		X"00",X"00",X"06",X"00",X"00",X"40",X"AE",X"2A",X"00",X"F8",X"FF",X"5F",X"C0",X"1D",X"00",X"80",
		X"E8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EF",X"7B",X"0F",X"40",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"FF",X"FF",X"FF",X"CF",X"01",X"00",X"80",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"0A",X"00",X"00",X"00",X"40",X"6F",X"85",X"00",X"00",X"00",X"EA",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"57",X"76",X"FF",X"FF",X"3B",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"F7",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"18",X"F8",X"FF",
		X"BF",X"F7",X"DD",X"01",X"0C",X"88",X"01",X"00",X"00",X"00",X"00",X"00",X"80",X"20",X"44",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"0E",X"FC",X"00",X"00",X"00",X"00",X"FE",X"FF",X"17",
		X"C0",X"C4",X"FF",X"FF",X"01",X"00",X"00",X"00",X"C8",X"C7",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"FF",X"07",X"40",X"0F",X"04",X"00",X"00",X"C0",X"07",X"10",X"00",X"C0",X"FF",X"FF",X"FF",
		X"BC",X"FF",X"FF",X"1F",X"07",X"02",X"00",X"00",X"00",X"80",X"FF",X"FF",X"FB",X"00",X"00",X"F0",
		X"FF",X"F3",X"01",X"00",X"FE",X"01",X"00",X"00",X"E8",X"0B",X"FF",X"FF",X"FF",X"33",X"00",X"FE",
		X"00",X"00",X"00",X"00",X"F0",X"FF",X"7F",X"00",X"78",X"FC",X"03",X"80",X"FF",X"F3",X"5F",X"89",
		X"3E",X"30",X"06",X"00",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"FF",X"1F",X"00",X"00",X"00",
		X"F8",X"01",X"00",X"00",X"10",X"FE",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"FF",X"07",X"00",X"80",
		X"01",X"00",X"00",X"78",X"7C",X"BE",X"F6",X"FF",X"FF",X"FF",X"7F",X"8C",X"FF",X"3F",X"00",X"00",
		X"00",X"18",X"00",X"00",X"00",X"F8",X"FF",X"FF",X"FF",X"2F",X"E0",X"FF",X"FF",X"FF",X"0D",X"00",
		X"00",X"00",X"00",X"F4",X"FF",X"7F",X"F8",X"FF",X"7F",X"00",X"00",X"B5",X"FD",X"0C",X"00",X"11",
		X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"80",X"A0",X"FB",X"00",X"00",X"00",X"00",X"1C",
		X"C3",X"01",X"00",X"F8",X"FF",X"FF",X"BF",X"12",X"FC",X"E3",X"3F",X"1F",X"C0",X"FF",X"01",X"00",
		X"00",X"FE",X"00",X"00",X"E0",X"7F",X"BF",X"00",X"A0",X"DD",X"1F",X"CF",X"FF",X"7F",X"01",X"3C",
		X"C0",X"07",X"70",X"80",X"7F",X"F0",X"38",X"1C",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"7F",X"FC",
		X"FF",X"7F",X"40",X"18",X"00",X"00",X"B8",X"00",X"00",X"FA",X"FF",X"CF",X"FF",X"E7",X"FF",X"FF",
		X"3F",X"00",X"00",X"70",X"06",X"E7",X"FF",X"FF",X"F1",X"03",X"00",X"00",X"D0",X"FF",X"FF",X"B9",
		X"FF",X"FF",X"9F",X"03",X"00",X"00",X"00",X"00",X"20",X"F0",X"FF",X"FF",X"FF",X"3F",X"3E",X"00",
		X"8C",X"33",X"00",X"F9",X"FF",X"FF",X"EF",X"C7",X"7F",X"38",X"38",X"80",X"21",X"A0",X"0A",X"08",
		X"00",X"00",X"00",X"F8",X"01",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F9",X"FF",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"00",X"48",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"80",X"EF",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",
		X"00",X"00",X"20",X"F0",X"FF",X"7F",X"70",X"00",X"00",X"E0",X"01",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"3F",X"FF",X"BF",X"01",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"FC",X"F7",X"9F",
		X"FF",X"E1",X"F9",X"3F",X"3F",X"00",X"00",X"00",X"00",X"FC",X"FF",X"7F",X"00",X"00",X"80",X"DE",
		X"1F",X"7F",X"BE",X"FF",X"FF",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"FE",X"FF",X"FF",X"FF",
		X"7F",X"05",X"00",X"00",X"00",X"00",X"40",X"2D",X"09",X"04",X"51",X"ED",X"FF",X"FF",X"FF",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"2F",X"FF",X"7F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"FE",X"FF",X"F3",X"F8",X"81",X"E3",X"4F",X"DA",X"F1",X"FF",X"FF",X"FF",X"FF",X"87",X"FF",X"07",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"20",X"E4",X"3F",X"00",X"FF",X"FF",X"FF",X"FF",X"00",
		X"F0",X"FF",X"FF",X"7F",X"B8",X"03",X"00",X"F0",X"FF",X"0F",X"00",X"00",X"80",X"E1",X"FF",X"07",
		X"00",X"80",X"FE",X"FF",X"F1",X"FD",X"FF",X"F9",X"FF",X"05",X"00",X"00",X"20",X"00",X"00",X"00",
		X"F0",X"FF",X"FF",X"FF",X"FF",X"87",X"07",X"6C",X"23",X"00",X"00",X"40",X"00",X"00",X"00",X"D8",
		X"FF",X"FF",X"7F",X"7F",X"FF",X"FF",X"03",X"00",X"00",X"F8",X"FF",X"CF",X"01",X"00",X"00",X"00",
		X"20",X"3C",X"DE",X"7F",X"FC",X"FF",X"03",X"E0",X"FF",X"FD",X"0F",X"00",X"00",X"FE",X"FF",X"03",
		X"00",X"00",X"A8",X"37",X"FF",X"E3",X"F8",X"83",X"B6",X"22",X"E0",X"00",X"00",X"00",X"C0",X"FF",
		X"FF",X"01",X"C0",X"FF",X"FF",X"38",X"00",X"C0",X"FF",X"FF",X"1E",X"00",X"00",X"00",X"00",X"E8",
		X"DF",X"DF",X"7F",X"FF",X"40",X"6F",X"45",X"E0",X"03",X"00",X"00",X"FC",X"FF",X"FF",X"FF",X"EF",
		X"8F",X"CF",X"7F",X"00",X"60",X"2B",X"A4",X"03",X"00",X"00",X"00",X"F8",X"F9",X"FF",X"FF",X"FF",
		X"FF",X"02",X"00",X"03",X"00",X"00",X"F0",X"FF",X"FF",X"FF",X"FF",X"BF",X"05",X"00",X"00",X"D0",
		X"AF",X"22",X"20",X"1E",X"00",X"00",X"FF",X"FF",X"FF",X"5F",X"D2",X"FE",X"FF",X"FF",X"FF",X"DF",
		X"81",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"05",X"78",X"00",X"00",X"00",X"F8",X"7D",X"57",X"55",X"A9",X"EC",X"3F",X"00",X"00",X"F8",
		X"FF",X"FF",X"FF",X"FD",X"1B",X"00",X"7F",X"DB",X"03",X"00",X"00",X"E8",X"00",X"00",X"C0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"02",X"00",X"80",X"DE",X"85",X"04",X"80",X"03",X"00",X"00",
		X"06",X"FE",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"40",X"CA",X"AA",X"55",X"95",X"84",X"00",X"00",
		X"FE",X"FF",X"01",X"00",X"00",X"FE",X"FF",X"3B",X"FE",X"7F",X"00",X"00",X"FC",X"FF",X"7F",X"00",
		X"1E",X"0F",X"00",X"00",X"3C",X"40",X"88",X"94",X"2A",X"FC",X"83",X"FF",X"F1",X"FF",X"FF",X"FF",
		X"EF",X"BA",X"1F",X"FC",X"7F",X"DB",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"02",X"00",X"00",X"1A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"11",X"02",
		X"F8",X"00",X"00",X"F0",X"FF",X"0F",X"1C",X"00",X"00",X"F8",X"FF",X"FF",X"00",X"00",X"70",X"E0",
		X"97",X"54",X"BD",X"FF",X"B7",X"FC",X"F8",X"FF",X"FF",X"4D",X"1C",X"08",X"00",X"F0",X"FF",X"DF",
		X"FF",X"7F",X"FE",X"FF",X"03",X"00",X"2A",X"0D",X"00",X"00",X"00",X"00",X"FE",X"FF",X"75",X"17",
		X"FE",X"FF",X"FF",X"FF",X"03",X"00",X"1F",X"40",X"F0",X"FF",X"3F",X"F0",X"01",X"FF",X"07",X"00",
		X"80",X"07",X"00",X"00",X"F8",X"1F",X"C0",X"FF",X"07",X"C0",X"FF",X"0F",X"00",X"08",X"F8",X"FF",
		X"5F",X"81",X"FF",X"9F",X"6F",X"A9",X"07",X"00",X"00",X"00",X"FE",X"FF",X"0F",X"00",X"C0",X"FF",
		X"03",X"30",X"FE",X"0D",X"DB",X"D6",X"1F",X"00",X"00",X"FF",X"FF",X"5F",X"DB",X"7B",X"83",X"FF",
		X"FF",X"07",X"00",X"20",X"00",X"FE",X"FF",X"0F",X"00",X"00",X"90",X"EE",X"FF",X"FF",X"1F",X"FF",
		X"FF",X"40",X"00",X"12",X"02",X"39",X"00",X"00",X"40",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"57",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"23",X"00",X"80",
		X"12",X"00",X"00",X"00",X"00",X"40",X"ED",X"FF",X"FF",X"1B",X"FD",X"FF",X"FF",X"FF",X"FF",X"7F",
		X"4B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E4",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"95",X"6A",X"FF",X"FF",X"FF",X"FF",X"3B",X"C0",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F5",X"FF",X"FF",X"FF",X"DF",X"F8",X"FF",X"FF",X"FF",X"7F",X"93",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"D0",X"B6",X"75",X"7D",X"00",X"A8",X"FF",X"FF",X"FF",X"FF",X"9F",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"F8",X"17",X"F8",X"FD",X"FF",X"DF",X"01",X"08",X"E0",
		X"E7",X"FF",X"FF",X"07",X"00",X"01",X"FC",X"FF",X"E3",X"08",X"81",X"10",X"22",X"00",X"B0",X"7F",
		X"00",X"18",X"01",X"00",X"DE",X"83",X"FF",X"FF",X"FF",X"FF",X"01",X"80",X"D4",X"DE",X"FF",X"FF",
		X"FF",X"6F",X"F0",X"FF",X"4A",X"00",X"00",X"02",X"00",X"01",X"80",X"FA",X"F9",X"FF",X"FF",X"FF",
		X"FF",X"01",X"00",X"00",X"00",X"3E",X"01",X"E8",X"B7",X"AA",X"06",X"00",X"00",X"00",X"B4",X"8B",
		X"FF",X"BF",X"FF",X"7F",X"13",X"C2",X"01",X"00",X"00",X"00",X"D4",X"F7",X"E3",X"FF",X"FF",X"07",
		X"00",X"00",X"00",X"FA",X"03",X"E0",X"FE",X"01",X"F8",X"81",X"53",X"6D",X"5F",X"9E",X"FF",X"FF",
		X"FF",X"0A",X"C0",X"01",X"00",X"00",X"40",X"DD",X"FF",X"FF",X"1D",X"FE",X"1F",X"88",X"58",X"1B",
		X"02",X"01",X"92",X"18",X"00",X"A0",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"5F",X"00",X"40",X"00",
		X"00",X"00",X"00",X"F5",X"FF",X"FF",X"EB",X"FF",X"FC",X"83",X"03",X"A0",X"D0",X"B1",X"AA",X"03",
		X"A4",X"F2",X"03",X"40",X"F8",X"FF",X"FF",X"F7",X"FF",X"E7",X"5F",X"41",X"00",X"40",X"7B",X"00",
		X"00",X"00",X"00",X"CC",X"1F",X"FF",X"FF",X"43",X"FF",X"DF",X"7F",X"00",X"DC",X"FF",X"0F",X"20",
		X"A4",X"6A",X"ED",X"B6",X"56",X"55",X"00",X"B0",X"AB",X"68",X"00",X"30",X"00",X"00",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"01",X"00",X"00",X"F5",X"01",X"00",X"00",X"D9",X"07",
		X"00",X"88",X"F0",X"FF",X"FF",X"3B",X"FF",X"FF",X"FF",X"1F",X"00",X"00",X"00",X"F0",X"5F",X"C1",
		X"FF",X"8F",X"40",X"66",X"FC",X"5A",X"15",X"A4",X"03",X"00",X"80",X"EC",X"BD",X"FC",X"FF",X"FF",
		X"99",X"04",X"00",X"09",X"00",X"00",X"00",X"ED",X"7D",X"F1",X"FF",X"1F",X"1E",X"C0",X"1E",X"00",
		X"D5",X"00",X"00",X"00",X"D2",X"DD",X"95",X"FF",X"FF",X"FF",X"5B",X"1F",X"80",X"00",X"00",X"00",
		X"FD",X"7C",X"3E",X"F8",X"FF",X"FF",X"0B",X"00",X"C0",X"4F",X"22",X"89",X"C3",X"FF",X"FF",X"8F",
		X"F1",X"00",X"00",X"A0",X"FF",X"FF",X"4B",X"44",X"24",X"7F",X"CB",X"A9",X"02",X"FF",X"FF",X"03",
		X"00",X"80",X"0E",X"FE",X"F1",X"23",X"24",X"25",X"FC",X"FF",X"FF",X"0B",X"38",X"10",X"22",X"E0",
		X"FF",X"FF",X"0F",X"01",X"20",X"92",X"AA",X"E0",X"FF",X"FF",X"B5",X"07",X"00",X"00",X"A6",X"DA",
		X"7D",X"FF",X"BD",X"7E",X"FC",X"FF",X"AA",X"06",X"80",X"00",X"1C",X"40",X"94",X"ED",X"AE",X"FF",
		X"FF",X"8A",X"FF",X"BF",X"D5",X"01",X"00",X"00",X"80",X"D4",X"56",X"FC",X"FF",X"FF",X"BB",X"96",
		X"52",X"1D",X"00",X"20",X"AA",X"DD",X"2F",X"FF",X"F3",X"FF",X"8F",X"55",X"2E",X"00",X"00",X"00",
		X"90",X"5A",X"EF",X"7D",X"37",X"F6",X"FF",X"DF",X"55",X"75",X"00",X"00",X"20",X"6B",X"37",X"FE",
		X"FF",X"FF",X"5F",X"00",X"00",X"88",X"01",X"FF",X"FF",X"12",X"00",X"C0",X"E3",X"7F",X"89",X"08",
		X"D1",X"FF",X"FF",X"2F",X"02",X"C0",X"FD",X"9F",X"24",X"F0",X"AF",X"AA",X"82",X"FF",X"BF",X"7B",
		X"00",X"00",X"C8",X"F0",X"E1",X"FD",X"0F",X"41",X"49",X"55",X"DB",X"DD",X"BB",X"BB",X"BA",X"CB",
		X"C1",X"85",X"1F",X"C0",X"03",X"80",X"48",X"C0",X"FF",X"FF",X"8F",X"07",X"DC",X"3F",X"27",X"C2",
		X"F1",X"3F",X"49",X"22",X"F0",X"7F",X"22",X"80",X"7F",X"02",X"E0",X"6E",X"AB",X"2A",X"23",X"AA",
		X"C3",X"83",X"54",X"FB",X"9E",X"FF",X"FF",X"FF",X"0F",X"80",X"02",X"42",X"10",X"12",X"A5",X"52",
		X"55",X"55",X"F8",X"55",X"29",X"E0",X"FF",X"BF",X"00",X"70",X"E6",X"7E",X"FC",X"DE",X"DB",X"B6",
		X"B5",X"5A",X"3F",X"00",X"22",X"59",X"6D",X"B7",X"EB",X"AA",X"4C",X"E0",X"00",X"02",X"18",X"08",
		X"6E",X"D7",X"F5",X"F0",X"03",X"C0",X"FF",X"5F",X"FF",X"F7",X"96",X"FF",X"FF",X"0D",X"AA",X"5A",
		X"00",X"00",X"00",X"80",X"48",X"BA",X"AA",X"5C",X"6B",X"B5",X"5A",X"6B",X"35",X"F1",X"FF",X"6F",
		X"D7",X"AA",X"1F",X"80",X"A8",X"DA",X"F2",X"FF",X"7F",X"FF",X"6F",X"15",X"11",X"0A",X"00",X"00",
		X"14",X"68",X"B5",X"54",X"AD",X"DB",X"DD",X"2E",X"FC",X"DF",X"D8",X"DD",X"76",X"00",X"00",X"4A",
		X"AD",X"FB",X"8E",X"FF",X"FF",X"07",X"FE",X"C0",X"AA",X"24",X"C9",X"01",X"20",X"3B",X"80",X"A4",
		X"DA",X"EE",X"FB",X"DE",X"DD",X"5A",X"12",X"7E",X"5B",X"27",X"00",X"00",X"D0",X"F7",X"BD",X"EF",
		X"74",X"DF",X"BC",X"D4",X"B6",X"7B",X"B7",X"F1",X"FF",X"0F",X"00",X"00",X"00",X"90",X"B6",X"1C",
		X"00",X"50",X"BB",X"9F",X"93",X"A4",X"EA",X"6E",X"7D",X"FF",X"FF",X"57",X"29",X"25",X"09",X"F8",
		X"7F",X"02",X"08",X"FA",X"00",X"3B",X"56",X"EB",X"38",X"20",X"88",X"BF",X"B6",X"DD",X"AE",X"F1",
		X"FF",X"5F",X"6D",X"10",X"18",X"00",X"0C",X"8E",X"53",X"C2",X"3F",X"8F",X"FF",X"6F",X"22",X"91",
		X"54",X"AA",X"AA",X"82",X"7F",X"FC",X"0F",X"02",X"D0",X"EE",X"E1",X"11",X"91",X"AA",X"8A",X"FE",
		X"FD",X"FF",X"22",X"84",X"80",X"BB",X"B7",X"D5",X"0E",X"08",X"10",X"E2",X"AA",X"B5",X"BB",X"DB",
		X"6D",X"F5",X"AA",X"29",X"C1",X"93",X"10",X"F0",X"83",X"EB",X"5A",X"AD",X"DA",X"07",X"80",X"C2",
		X"FF",X"E7",X"7F",X"29",X"A5",X"2A",X"C1",X"4F",X"12",X"40",X"5B",X"AD",X"03",X"00",X"80",X"92",
		X"6A",X"BB",X"ED",X"FE",X"FF",X"FF",X"6C",X"1F",X"80",X"87",X"D6",X"D6",X"DA",X"16",X"88",X"A8",
		X"54",X"EB",X"B6",X"5A",X"95",X"70",X"0E",X"00",X"F5",X"01",X"04",X"F8",X"90",X"A4",X"E0",X"FF",
		X"FF",X"0A",X"FF",X"7F",X"D7",X"1D",X"81",X"60",X"BB",X"FB",X"10",X"88",X"22",X"A9",X"12",X"5E",
		X"09",X"B7",X"5B",X"95",X"D0",X"00",X"0C",X"20",X"A9",X"DD",X"FF",X"77",X"FE",X"FF",X"7F",X"1F",
		X"1C",X"00",X"3C",X"A0",X"F6",X"01",X"AE",X"23",X"A5",X"AA",X"AA",X"E2",X"DF",X"7F",X"48",X"04",
		X"41",X"A2",X"94",X"AA",X"D6",X"DA",X"E2",X"FF",X"2A",X"D8",X"DB",X"B5",X"AA",X"92",X"7A",X"00",
		X"22",X"D5",X"EE",X"7D",X"EB",X"FF",X"DF",X"AA",X"04",X"11",X"01",X"00",X"2C",X"48",X"AA",X"DA",
		X"DE",X"F7",X"DD",X"ED",X"8A",X"3F",X"AE",X"35",X"1D",X"00",X"70",X"90",X"28",X"C5",X"FF",X"FF",
		X"AB",X"A4",X"E0",X"4F",X"C2",X"EE",X"76",X"80",X"40",X"08",X"F6",X"4B",X"49",X"A9",X"2A",X"FC",
		X"57",X"AB",X"AA",X"E2",X"D5",X"AA",X"8A",X"FB",X"6E",X"5B",X"55",X"D5",X"03",X"00",X"E0",X"DE",
		X"DF",X"F7",X"1E",X"03",X"A0",X"E3",X"03",X"D5",X"44",X"92",X"94",X"4A",X"55",X"15",X"FE",X"57",
		X"25",X"B2",X"54",X"AA",X"AA",X"7E",X"DB",X"55",X"FB",X"7F",X"95",X"12",X"7B",X"63",X"DB",X"4A",
		X"D1",X"81",X"01",X"00",X"A6",X"AA",X"84",X"FF",X"FF",X"E5",X"20",X"20",X"44",X"52",X"65",X"E2",
		X"BF",X"BB",X"D5",X"AA",X"54",X"4A",X"F5",X"41",X"52",X"DD",X"EF",X"DF",X"F7",X"6E",X"AB",X"F8",
		X"21",X"08",X"80",X"0E",X"06",X"92",X"2A",X"00",X"58",X"B1",X"5F",X"AB",X"6D",X"B7",X"FA",X"7F",
		X"AF",X"AA",X"28",X"EF",X"F1",X"80",X"81",X"40",X"C0",X"FE",X"24",X"DC",X"6D",X"DB",X"17",X"88",
		X"24",X"F2",X"DF",X"AA",X"5A",X"F8",X"BE",X"D7",X"07",X"10",X"40",X"1F",X"D8",X"4E",X"92",X"94",
		X"AA",X"6A",X"6D",X"6B",X"6B",X"55",X"F0",X"CF",X"56",X"55",X"04",X"A8",X"06",X"82",X"54",X"E9",
		X"EF",X"BE",X"BB",X"FC",X"CB",X"27",X"91",X"42",X"04",X"B4",X"56",X"55",X"07",X"03",X"40",X"BB",
		X"F7",X"7E",X"2A",X"55",X"6B",X"DB",X"16",X"FF",X"BF",X"8B",X"80",X"00",X"2E",X"0A",X"43",X"1C",
		X"BC",X"5C",X"4A",X"5A",X"A9",X"EA",X"AA",X"3C",X"FF",X"DE",X"0F",X"81",X"DA",X"86",X"48",X"A9",
		X"AA",X"F8",X"FB",X"2A",X"E1",X"1F",X"45",X"A8",X"24",X"89",X"F0",X"1E",X"B7",X"8E",X"07",X"38",
		X"70",X"A7",X"14",X"BF",X"CA",X"EF",X"77",X"1F",X"44",X"6D",X"A0",X"2A",X"AD",X"20",X"A2",X"52",
		X"B5",X"D6",X"D6",X"56",X"15",X"7E",X"3F",X"82",X"C0",X"3C",X"A8",X"5B",X"12",X"A9",X"AA",X"76",
		X"BB",X"DB",X"6D",X"2D",X"FE",X"6D",X"55",X"0A",X"20",X"05",X"1A",X"20",X"52",X"15",X"FF",X"7E",
		X"AD",X"E8",X"BD",X"6D",X"07",X"02",X"0C",X"F6",X"48",X"49",X"89",X"FB",X"FB",X"12",X"6E",X"FB",
		X"22",X"9C",X"25",X"A5",X"64",X"F9",X"DE",X"B6",X"6A",X"05",X"80",X"90",X"94",X"AA",X"5A",X"AD",
		X"C5",X"F7",X"1E",X"78",X"88",X"08",X"3F",X"E2",X"14",X"F4",X"BE",X"8B",X"27",X"1E",X"AE",X"AB",
		X"AA",X"B8",X"FC",X"B9",X"D5",X"4A",X"0D",X"40",X"90",X"08",X"F7",X"4F",X"15",X"71",X"9F",X"C0",
		X"5A",X"AB",X"D5",X"82",X"10",X"4D",X"55",X"D5",X"6F",X"AB",X"DE",X"F7",X"2B",X"84",X"88",X"92",
		X"A4",X"5A",X"55",X"55",X"DC",X"6F",X"5B",X"75",X"80",X"20",X"92",X"AA",X"DA",X"EE",X"76",X"E5",
		X"EF",X"DB",X"AA",X"24",X"22",X"32",X"00",X"44",X"D2",X"FA",X"6D",X"B7",X"AD",X"F1",X"7B",X"5B",
		X"55",X"0A",X"00",X"00",X"DA",X"BA",X"27",X"29",X"F1",X"BD",X"FB",X"A4",X"94",X"54",X"C9",X"93",
		X"47",X"6D",X"77",X"42",X"88",X"24",X"C9",X"53",X"55",X"55",X"F4",X"E7",X"87",X"B5",X"1E",X"40",
		X"73",X"82",X"DD",X"A7",X"AA",X"14",X"7E",X"EF",X"97",X"50",X"AC",X"AA",X"A2",X"10",X"22",X"A5",
		X"AA",X"5A",X"2B",X"FE",X"FB",X"52",X"82",X"7A",X"E8",X"38",X"4A",X"70",X"7F",X"B8",X"2E",X"71",
		X"78",X"89",X"17",X"4F",X"95",X"AA",X"A2",X"BA",X"6D",X"D5",X"02",X"86",X"10",X"52",X"AA",X"52",
		X"FF",X"D6",X"D5",X"6A",X"55",X"C5",X"F7",X"CB",X"08",X"31",X"51",X"69",X"F0",X"AF",X"4A",X"A6",
		X"87",X"B7",X"6B",X"55",X"55",X"15",X"30",X"45",X"92",X"54",X"55",X"DF",X"8A",X"EF",X"D9",X"6A",
		X"01",X"81",X"88",X"A4",X"AA",X"5D",X"75",X"B5",X"AE",X"FC",X"E9",X"15",X"7E",X"A9",X"25",X"A5",
		X"AA",X"12",X"F7",X"7D",X"C0",X"1E",X"54",X"3D",X"04",X"AC",X"76",X"4A",X"4A",X"55",X"55",X"C5",
		X"EF",X"97",X"12",X"11",X"0B",X"6B",X"AB",X"AA",X"AA",X"54",X"07",X"81",X"FB",X"AA",X"B5",X"ED",
		X"B6",X"7B",X"AD",X"56",X"55",X"22",X"02",X"55",X"55",X"12",X"05",X"12",X"82",X"48",X"69",X"DD",
		X"7B",X"EF",X"DD",X"55",X"FF",X"D8",X"1E",X"41",X"98",X"80",X"56",X"2F",X"92",X"A4",X"4A",X"75",
		X"EF",X"B9",X"57",X"04",X"AD",X"AD",X"CB",X"D0",X"0B",X"E1",X"54",X"EC",X"6D",X"DB",X"AA",X"75",
		X"40",X"55",X"25",X"22",X"AA",X"AA",X"6A",X"55",X"77",X"BC",X"77",X"53",X"10",X"A2",X"5A",X"A5",
		X"54",X"AA",X"AA",X"F5",X"5A",X"77",X"AB",X"56",X"15",X"CA",X"8B",X"0A",X"FC",X"82",X"D5",X"09",
		X"55",X"1D",X"49",X"14",X"BD",X"AA",X"E5",X"FE",X"FE",X"14",X"C1",X"03",X"AB",X"56",X"75",X"81",
		X"22",X"55",X"A1",X"F7",X"6E",X"5B",X"57",X"42",X"92",X"52",X"E8",X"DE",X"6D",X"5D",X"12",X"44",
		X"52",X"92",X"AB",X"AA",X"8A",X"BF",X"2E",X"A4",X"EA",X"22",X"49",X"A9",X"AA",X"6A",X"B7",X"6D",
		X"AD",X"15",X"7E",X"B7",X"3D",X"02",X"60",X"0B",X"B6",X"F6",X"29",X"44",X"FB",X"84",X"DD",X"B6",
		X"A7",X"02",X"27",X"29",X"B2",X"67",X"8A",X"A7",X"17",X"12",X"58",X"ED",X"51",X"8A",X"26",X"5D",
		X"AD",X"BA",X"5A",X"6B",X"2D",X"BD",X"9F",X"4A",X"24",X"A1",X"7D",X"45",X"08",X"D6",X"5A",X"8F",
		X"44",X"49",X"8A",X"5C",X"7F",X"55",X"55",X"91",X"8F",X"3F",X"25",X"49",X"8A",X"A2",X"FB",X"A9",
		X"48",X"58",X"BB",X"AD",X"56",X"55",X"95",X"8E",X"7A",X"94",X"A4",X"AA",X"75",X"B7",X"6D",X"AB",
		X"AA",X"A0",X"3E",X"10",X"58",X"10",X"61",X"89",X"B8",X"25",X"FC",X"55",X"15",X"FF",X"E2",X"ED",
		X"6A",X"6D",X"93",X"28",X"29",X"F1",X"F1",X"4B",X"74",X"57",X"11",X"49",X"54",X"4A",X"95",X"AA",
		X"2A",X"E1",X"DE",X"ED",X"12",X"92",X"E0",X"AB",X"DC",X"AD",X"CA",X"7B",X"B7",X"56",X"55",X"87",
		X"A0",X"AA",X"0C",X"49",X"4A",X"55",X"D5",X"AA",X"AA",X"2A",X"D8",X"BA",X"4A",X"12",X"49",X"51",
		X"80",X"A4",X"6A",X"F7",X"FB",X"6E",X"FF",X"5F",X"55",X"C5",X"B6",X"AC",X"10",X"11",X"29",X"32",
		X"9D",X"12",X"ED",X"54",X"A2",X"2F",X"F2",X"55",X"52",X"2A",X"C5",X"4F",X"8B",X"5B",X"AD",X"AA",
		X"52",X"A9",X"54",X"A5",X"6A",X"3D",X"E8",X"C7",X"56",X"55",X"AB",X"B5",X"5A",X"55",X"A5",X"A4",
		X"48",X"12",X"81",X"6A",X"B5",X"AA",X"54",X"AA",X"85",X"A4",X"6A",X"7F",X"EF",X"B6",X"FF",X"BB",
		X"27",X"30",X"AA",X"41",X"91",X"48",X"52",X"2A",X"55",X"D2",X"E5",X"ED",X"93",X"48",X"95",X"F0",
		X"2B",X"5F",X"15",X"DE",X"6E",X"5B",X"AB",X"D6",X"60",X"D5",X"A1",X"94",X"4A",X"4E",X"5F",X"55",
		X"78",X"61",X"55",X"55",X"11",X"84",X"88",X"52",X"55",X"B5",X"B6",X"ED",X"B6",X"FA",X"DA",X"AA",
		X"AA",X"E8",X"6E",X"D5",X"EA",X"40",X"14",X"AA",X"54",X"55",X"DF",X"6A",X"E3",X"6D",X"DB",X"05",
		X"94",X"41",X"8B",X"D0",X"E2",X"54",X"AA",X"8A",X"DF",X"57",X"55",X"E1",X"B6",X"D6",X"AA",X"8A",
		X"52",X"C5",X"C0",X"4A",X"55",X"55",X"D5",X"BF",X"4E",X"57",X"9A",X"92",X"92",X"24",X"49",X"52",
		X"D4",X"52",X"A5",X"4A",X"55",X"B8",X"EF",X"6E",X"A7",X"04",X"2D",X"FA",X"AA",X"6A",X"55",X"7C",
		X"77",X"73",X"85",X"41",X"05",X"27",X"89",X"5D",X"4A",X"B2",X"7D",X"4A",X"C4",X"6A",X"7B",X"09",
		X"D5",X"AA",X"AE",X"9D",X"48",X"55",X"55",X"B7",X"BA",X"BE",X"4E",X"55",X"11",X"AD",X"44",X"91",
		X"B8",X"4C",X"4C",X"D4",X"A2",X"F6",X"B0",X"AC",X"6E",X"6A",X"55",X"76",X"B5",X"AA",X"B6",X"02",
		X"52",X"12",X"A1",X"52",X"D5",X"BF",X"50",X"41",X"D3",X"AF",X"AE",X"05",X"62",X"95",X"D6",X"62",
		X"A3",X"15",X"A5",X"7A",X"D2",X"57",X"58",X"54",X"7C",X"45",X"AF",X"E8",X"9F",X"6A",X"B9",X"40",
		X"4B",X"08",X"7D",X"A0",X"F2",X"87",X"F8",X"7E",X"40",X"BF",X"92",X"C2",X"07",X"A9",X"7F",X"D6",
		X"D2",X"A0",X"74",X"A9",X"06",X"B5",X"E7",X"E0",X"D4",X"71",X"7C",X"AA",X"D5",X"9A",X"1C",X"B8",
		X"3A",X"9A",X"52",X"AF",X"54",X"85",X"DA",X"90",X"D4",X"4B",X"0A",X"C7",X"AF",X"22",X"34",X"29",
		X"A7",X"EA",X"6B",X"7D",X"41",X"DD",X"A2",X"4A",X"5D",X"F4",X"76",X"29",X"6E",X"80",X"97",X"CA",
		X"49",X"5C",X"75",X"11",X"69",X"CF",X"13",X"9A",X"1E",X"B4",X"A2",X"55",X"B9",X"DA",X"20",X"F5",
		X"A7",X"60",X"D7",X"1A",X"6E",X"A7",X"85",X"A3",X"E4",X"A2",X"5A",X"D8",X"8E",X"EA",X"A5",X"9B",
		X"74",X"D5",X"35",X"C0",X"AA",X"25",X"BC",X"2A",X"DE",X"A6",X"1D",X"1B",X"F2",X"42",X"EA",X"A5",
		X"A3",X"E2",X"7A",X"21",X"B1",X"F6",X"29",X"3C",X"CA",X"75",X"85",X"3E",X"A8",X"3C",X"69",X"A8",
		X"FD",X"16",X"D5",X"63",X"A1",X"74",X"14",X"BA",X"AE",X"07",X"56",X"C3",X"50",X"35",X"DD",X"45",
		X"7A",X"59",X"9D",X"03",X"F3",X"C2",X"2B",X"C5",X"57",X"33",X"50",X"FF",X"01",X"4C",X"7E",X"34",
		X"4A",X"AB",X"83",X"C7",X"34",X"F8",X"F1",X"50",X"B1",X"0E",X"53",X"7D",X"5C",X"CB",X"82",X"0F",
		X"BC",X"D0",X"F0",X"87",X"BB",X"F0",X"E1",X"83",X"53",X"1E",X"DD",X"B4",X"0A",X"16",X"6E",X"87",
		X"BE",X"86",X"73",X"1D",X"F0",X"0B",X"6C",X"29",X"74",X"85",X"AF",X"83",X"EA",X"A5",X"C1",X"52",
		X"27",X"AC",X"07",X"5F",X"A5",X"B7",X"C4",X"E0",X"EB",X"01",X"F8",X"3F",X"C0",X"1F",X"38",X"FD",
		X"00",X"1F",X"F0",X"EA",X"02",X"3F",X"E0",X"6B",X"01",X"7F",X"E8",X"43",X"D1",X"F3",X"54",X"56",
		X"54",X"BD",X"A0",X"1E",X"97",X"28",X"E5",X"AA",X"7A",X"5D",X"0B",X"A2",X"F5",X"14",X"5E",X"AA",
		X"6F",X"3C",X"90",X"B5",X"25",X"21",X"A5",X"9B",X"AF",X"06",X"9D",X"E6",X"FA",X"2A",X"AD",X"E8",
		X"93",X"5C",X"91",X"00",X"50",X"25",X"24",X"AF",X"3F",X"FC",X"FF",X"F5",X"F0",X"53",X"79",X"E0",
		X"05",X"C2",X"81",X"4E",X"4D",X"20",X"6B",X"79",X"01",X"6E",X"E0",X"87",X"F9",X"F8",X"D4",X"3B",
		X"F6",X"16",X"63",X"67",X"7B",X"E0",X"F8",X"30",X"06",X"47",X"51",X"74",X"E1",X"8E",X"A8",X"BD",
		X"54",X"F0",X"67",X"7C",X"E0",X"0F",X"FA",X"57",X"F0",X"A6",X"78",X"83",X"50",X"11",X"43",X"FC",
		X"50",X"EB",X"C2",X"C7",X"FF",X"06",X"58",X"FF",X"81",X"0E",X"AF",X"0A",X"C0",X"55",X"42",X"8B",
		X"82",X"FF",X"EB",X"7F",X"AD",X"EE",X"80",X"22",X"48",X"0D",X"C0",X"30",X"F8",X"82",X"45",X"12",
		X"3F",X"FC",X"DF",X"FF",X"7D",X"87",X"E3",X"EF",X"1F",X"BC",X"81",X"09",X"00",X"00",X"84",X"05",
		X"F4",X"DF",X"1F",X"1E",X"69",X"57",X"C9",X"55",X"24",X"B8",X"FC",X"41",X"FF",X"FF",X"07",X"2D",
		X"1D",X"70",X"78",X"80",X"70",X"01",X"6C",X"95",X"38",X"E9",X"7F",X"FD",X"FB",X"A0",X"3F",X"81",
		X"00",X"7E",X"23",X"EA",X"FB",X"4A",X"20",X"ED",X"0B",X"00",X"00",X"91",X"AA",X"BA",X"7D",X"FD",
		X"FF",X"87",X"FB",X"BF",X"BE",X"2A",X"31",X"50",X"06",X"40",X"1E",X"68",X"15",X"04",X"28",X"AA",
		X"F4",X"FF",X"FF",X"FF",X"E7",X"14",X"14",X"8E",X"94",X"4A",X"05",X"EA",X"06",X"00",X"00",X"07",
		X"EC",X"FF",X"FF",X"8F",X"80",X"88",X"88",X"04",X"BF",X"7F",X"FF",X"C8",X"43",X"3F",X"00",X"A0",
		X"7D",X"90",X"F5",X"C1",X"5A",X"3F",X"1E",X"21",X"48",X"AA",X"D6",X"5B",X"FC",X"F7",X"FF",X"1F",
		X"1C",X"1F",X"00",X"C0",X"03",X"6C",X"FF",X"01",X"80",X"04",X"F0",X"FB",X"EF",X"FD",X"27",X"00",
		X"84",X"24",X"6D",X"15",X"FE",X"FF",X"FF",X"7F",X"80",X"1F",X"40",X"FC",X"10",X"00",X"01",X"9C",
		X"FF",X"FF",X"C1",X"11",X"22",X"49",X"55",X"F0",X"E3",X"F7",X"DF",X"AD",X"9A",X"E4",X"03",X"00",
		X"00",X"90",X"AA",X"C2",X"FF",X"E9",X"FF",X"FF",X"07",X"E0",X"17",X"00",X"20",X"45",X"2A",X"95",
		X"3E",X"F8",X"F7",X"DD",X"ED",X"E1",X"B0",X"00",X"00",X"80",X"C0",X"37",X"7C",X"F8",X"FF",X"F9",
		X"C0",X"FF",X"04",X"F8",X"C1",X"20",X"91",X"04",X"FC",X"FD",X"BE",X"B7",X"5A",X"A5",X"3E",X"18",
		X"00",X"00",X"45",X"70",X"FA",X"FF",X"79",X"FD",X"DA",X"FD",X"07",X"40",X"5A",X"54",X"54",X"05",
		X"73",X"03",X"00",X"C3",X"FB",X"FF",X"2F",X"02",X"31",X"FF",X"17",X"60",X"FF",X"EB",X"0F",X"00",
		X"0E",X"94",X"2F",X"63",X"80",X"8D",X"43",X"22",X"09",X"F8",X"FF",X"FF",X"EF",X"77",X"01",X"C0",
		X"87",X"12",X"2E",X"10",X"3C",X"57",X"2D",X"83",X"FF",X"FF",X"17",X"22",X"11",X"00",X"FC",X"81",
		X"EE",X"DD",X"7F",X"08",X"E0",X"70",X"28",X"52",X"12",X"17",X"CD",X"FF",X"7F",X"F8",X"4F",X"48",
		X"54",X"5A",X"C0",X"F5",X"FB",X"3E",X"A8",X"BE",X"00",X"00",X"01",X"F8",X"80",X"FF",X"FF",X"83",
		X"BF",X"4F",X"01",X"C0",X"BF",X"50",X"02",X"FC",X"BF",X"F7",X"F3",X"05",X"00",X"85",X"87",X"C7",
		X"0F",X"05",X"11",X"96",X"82",X"FF",X"71",X"FF",X"7E",X"FF",X"02",X"00",X"00",X"FA",X"9F",X"83",
		X"7F",X"09",X"70",X"20",X"F4",X"FF",X"8B",X"84",X"44",X"E0",X"F1",X"FF",X"FD",X"EA",X"79",X"01",
		X"00",X"00",X"FF",X"87",X"28",X"61",X"B9",X"A5",X"E0",X"FF",X"7D",X"FF",X"07",X"00",X"00",X"D0",
		X"FD",X"AD",X"AE",X"6F",X"01",X"A2",X"EB",X"07",X"C0",X"3F",X"C1",X"70",X"AC",X"BA",X"C1",X"FF",
		X"A3",X"FF",X"8F",X"84",X"40",X"A8",X"B6",X"6B",X"7F",X"01",X"00",X"00",X"C0",X"97",X"CF",X"5B",
		X"F8",X"FF",X"3F",X"E0",X"0F",X"50",X"FF",X"03",X"D4",X"FE",X"70",X"02",X"A0",X"00",X"8E",X"BE",
		X"EF",X"1F",X"D4",X"FE",X"5F",X"00",X"00",X"01",X"B0",X"F7",X"FB",X"FF",X"69",X"00",X"AC",X"F1",
		X"41",X"20",X"80",X"B9",X"EF",X"6F",X"FF",X"BE",X"C0",X"F8",X"01",X"00",X"B8",X"04",X"FA",X"FF",
		X"FF",X"7F",X"01",X"10",X"44",X"4A",X"82",X"FB",X"FF",X"FB",X"07",X"F0",X"07",X"00",X"58",X"12",
		X"01",X"FE",X"0F",X"EF",X"FF",X"00",X"F7",X"2B",X"0F",X"01",X"20",X"49",X"49",X"F0",X"FF",X"FF",
		X"FF",X"04",X"C0",X"1F",X"1F",X"C8",X"A1",X"C0",X"02",X"F8",X"FE",X"FD",X"3D",X"0E",X"00",X"84",
		X"48",X"C0",X"FE",X"FF",X"7F",X"11",X"C0",X"FF",X"09",X"84",X"05",X"16",X"C2",X"FF",X"FF",X"01",
		X"0F",X"51",X"00",X"FF",X"5F",X"38",X"A0",X"B2",X"F7",X"FF",X"04",X"E0",X"23",X"F5",X"8F",X"00",
		X"42",X"12",X"AF",X"F8",X"F5",X"2F",X"BD",X"FF",X"FF",X"A8",X"00",X"80",X"75",X"C0",X"03",X"20",
		X"AA",X"BB",X"B5",X"ED",X"0F",X"18",X"F9",X"01",X"FF",X"01",X"FB",X"C1",X"CF",X"1F",X"78",X"00",
		X"F8",X"BF",X"1F",X"58",X"BB",X"07",X"02",X"80",X"00",X"C0",X"7F",X"F8",X"FD",X"7F",X"01",X"4A",
		X"25",X"A0",X"FE",X"EB",X"0F",X"7F",X"05",X"F0",X"0B",X"00",X"56",X"08",X"FF",X"E1",X"E7",X"7F",
		X"02",X"00",X"F8",X"7F",X"01",X"F5",X"07",X"7F",X"C0",X"A3",X"44",X"42",X"C0",X"FF",X"1F",X"F4",
		X"FE",X"05",X"C0",X"3F",X"80",X"7F",X"42",X"48",X"84",X"F3",X"D0",X"FF",X"BF",X"ED",X"54",X"CB",
		X"03",X"00",X"E0",X"17",X"04",X"F4",X"DF",X"87",X"EF",X"3D",X"01",X"F0",X"1F",X"DC",X"97",X"10",
		X"04",X"FE",X"4F",X"02",X"5D",X"49",X"C1",X"03",X"EF",X"DF",X"BB",X"54",X"D5",X"0B",X"00",X"00",
		X"7C",X"00",X"FF",X"7F",X"92",X"28",X"7E",X"E0",X"7F",X"EC",X"BF",X"77",X"43",X"D5",X"0B",X"08",
		X"00",X"80",X"04",X"F8",X"FF",X"7F",X"49",X"92",X"54",X"55",X"AD",X"E0",X"FE",X"DF",X"5B",X"BB",
		X"07",X"00",X"00",X"00",X"4C",X"FF",X"E3",X"FD",X"BF",X"80",X"2F",X"00",X"3F",X"1C",X"FC",X"E0",
		X"DD",X"F5",X"D3",X"FF",X"08",X"00",X"60",X"09",X"BC",X"FD",X"F8",X"0F",X"07",X"81",X"E0",X"FE",
		X"07",X"74",X"45",X"50",X"C0",X"FB",X"6F",X"FF",X"03",X"86",X"7E",X"22",X"00",X"F8",X"A8",X"60",
		X"D1",X"F9",X"FF",X"FF",X"FD",X"08",X"00",X"21",X"94",X"14",X"E8",X"FF",X"FF",X"9F",X"07",X"00",
		X"88",X"80",X"2F",X"78",X"FF",X"F5",X"FA",X"44",X"00",X"81",X"02",X"7E",X"FF",X"DF",X"FE",X"00",
		X"D4",X"FA",X"0B",X"20",X"44",X"92",X"05",X"FD",X"FF",X"FF",X"4C",X"A0",X"10",X"55",X"55",X"82",
		X"DC",X"FF",X"76",X"55",X"55",X"09",X"09",X"84",X"94",X"17",X"00",X"80",X"A4",X"F8",X"7F",X"FC",
		X"FF",X"15",X"FF",X"FF",X"AE",X"EA",X"E1",X"03",X"00",X"1C",X"0A",X"00",X"54",X"0A",X"E2",X"F7",
		X"3F",X"FB",X"1F",X"7E",X"02",X"21",X"A8",X"80",X"9F",X"BF",X"FF",X"81",X"97",X"80",X"90",X"A4",
		X"54",X"FC",X"44",X"BF",X"6D",X"FF",X"03",X"C2",X"3F",X"E0",X"50",X"F9",X"01",X"1C",X"21",X"02",
		X"F8",X"FF",X"DF",X"3F",X"6D",X"F5",X"07",X"80",X"5F",X"00",X"E0",X"7F",X"40",X"F8",X"BF",X"04",
		X"09",X"FE",X"8B",X"D0",X"EF",X"B6",X"ED",X"0F",X"10",X"10",X"80",X"10",X"21",X"F4",X"3F",X"3F",
		X"FA",X"FF",X"BB",X"01",X"C0",X"FD",X"E0",X"5A",X"00",X"9A",X"92",X"84",X"EE",X"6F",X"C2",X"FF",
		X"78",X"7F",X"F0",X"01",X"5A",X"3F",X"0B",X"07",X"00",X"20",X"5F",X"A1",X"4A",X"40",X"FF",X"FF",
		X"FF",X"CF",X"00",X"94",X"0F",X"F8",X"E1",X"80",X"FE",X"00",X"D5",X"9F",X"88",X"A4",X"14",X"1E",
		X"FF",X"FF",X"B7",X"3F",X"23",X"00",X"00",X"01",X"8F",X"FF",X"7F",X"11",X"22",X"2C",X"E0",X"FF",
		X"21",X"D6",X"FF",X"0B",X"00",X"FF",X"00",X"D8",X"AB",X"AB",X"A7",X"1E",X"1E",X"1C",X"40",X"7E",
		X"41",X"F7",X"FF",X"00",X"3E",X"FE",X"C0",X"9F",X"00",X"80",X"BF",X"0E",X"AB",X"7F",X"01",X"82",
		X"90",X"94",X"A0",X"FF",X"FF",X"17",X"12",X"80",X"BD",X"B7",X"DE",X"03",X"3E",X"20",X"60",X"00",
		X"FF",X"DF",X"AB",X"54",X"55",X"E0",X"FF",X"FF",X"03",X"57",X"3F",X"58",X"00",X"A1",X"0F",X"05",
		X"78",X"09",X"52",X"AA",X"55",X"BF",X"BD",X"E0",X"FF",X"FD",X"AF",X"00",X"04",X"80",X"B6",X"ED",
		X"FE",X"00",X"18",X"04",X"28",X"FE",X"C3",X"0F",X"EF",X"DF",X"AD",X"6A",X"D5",X"2F",X"40",X"80",
		X"90",X"38",X"7C",X"CF",X"FF",X"BF",X"7B",X"FD",X"80",X"00",X"D6",X"C0",X"21",X"00",X"02",X"FF",
		X"80",X"FF",X"2F",X"29",X"A5",X"28",X"F8",X"DF",X"EF",X"BF",X"07",X"00",X"00",X"3C",X"D0",X"DF",
		X"2F",X"42",X"80",X"D7",X"83",X"FE",X"7D",X"80",X"67",X"DF",X"1F",X"02",X"88",X"08",X"7C",X"55",
		X"75",X"83",X"FF",X"EF",X"40",X"FF",X"01",X"10",X"B4",X"FF",X"03",X"00",X"3F",X"50",X"BB",X"FD",
		X"0E",X"20",X"E0",X"07",X"F7",X"7D",X"77",X"D5",X"3A",X"80",X"B4",X"3D",X"42",X"00",X"1A",X"F0",
		X"FB",X"FF",X"FB",X"0B",X"00",X"21",X"00",X"DB",X"FF",X"FD",X"07",X"7C",X"40",X"00",X"78",X"41",
		X"FF",X"F7",X"E1",X"07",X"8F",X"00",X"5D",X"4A",X"5C",X"D5",X"C3",X"FD",X"7E",X"F0",X"F0",X"E1",
		X"D1",X"E3",X"0B",X"00",X"CC",X"03",X"1F",X"02",X"55",X"DC",X"E2",X"F8",X"FB",X"FF",X"17",X"02",
		X"28",X"F0",X"F0",X"FE",X"07",X"A6",X"55",X"AD",X"8D",X"09",X"3C",X"01",X"40",X"00",X"FA",X"FF",
		X"FF",X"1B",X"B1",X"04",X"5A",X"FD",X"7F",X"80",X"FA",X"87",X"D4",X"0F",X"01",X"90",X"D0",X"52",
		X"6E",X"FD",X"2D",X"F0",X"FF",X"58",X"81",X"D3",X"7D",X"E0",X"16",X"00",X"00",X"DD",X"2F",X"6D",
		X"AB",X"FA",X"03",X"0F",X"0A",X"AD",X"22",X"3A",X"FE",X"CF",X"92",X"FF",X"E7",X"C7",X"03",X"07",
		X"BC",X"07",X"C0",X"1E",X"20",X"EA",X"0C",X"56",X"05",X"18",X"7C",X"55",X"C1",X"FF",X"EF",X"07",
		X"FF",X"7F",X"C0",X"F1",X"F1",X"00",X"06",X"A4",X"FB",X"F1",X"42",X"90",X"00",X"EE",X"7F",X"FF",
		X"16",X"18",X"70",X"E9",X"F9",X"0B",X"08",X"0A",X"BE",X"52",X"55",X"55",X"81",X"F7",X"C7",X"7D",
		X"7D",X"10",X"A0",X"DA",X"B9",X"00",X"00",X"5B",X"E0",X"FD",X"4B",X"05",X"1F",X"FC",X"FF",X"5F",
		X"7D",X"0D",X"C0",X"59",X"00",X"CE",X"C3",X"07",X"3C",X"F0",X"E1",X"51",X"53",X"2A",X"FC",X"35",
		X"E8",X"FF",X"7F",X"00",X"7E",X"18",X"78",X"2B",X"00",X"01",X"0F",X"AE",X"FF",X"F6",X"F9",X"04",
		X"83",X"96",X"24",X"EC",X"7F",X"2D",X"5E",X"55",X"91",X"1E",X"1F",X"BE",X"EF",X"6A",X"15",X"84",
		X"7C",X"00",X"00",X"20",X"20",X"E9",X"FF",X"77",X"15",X"E4",X"B7",X"FF",X"7F",X"40",X"68",X"8F",
		X"05",X"90",X"8A",X"F4",X"10",X"F4",X"0F",X"F4",X"BF",X"EB",X"0F",X"00",X"F5",X"50",X"BD",X"A2",
		X"AD",X"E0",X"81",X"88",X"54",X"55",X"85",X"FF",X"C3",X"FF",X"FF",X"01",X"7E",X"01",X"45",X"95",
		X"20",X"09",X"F0",X"7E",X"DB",X"7F",X"20",X"00",X"FA",X"03",X"B4",X"7F",X"04",X"C8",X"A0",X"FF",
		X"FB",X"1F",X"70",X"F8",X"45",X"12",X"81",X"FF",X"A1",X"B7",X"3F",X"40",X"3E",X"04",X"90",X"F6",
		X"DE",X"EE",X"82",X"22",X"10",X"A5",X"68",X"FC",X"8B",X"FE",X"71",X"BF",X"EF",X"0F",X"3E",X"00",
		X"00",X"44",X"C2",X"2B",X"B6",X"FF",X"BE",X"BB",X"6D",X"1F",X"12",X"00",X"C0",X"87",X"81",X"FB",
		X"BF",X"40",X"7F",X"0E",X"8E",X"BF",X"A0",X"C0",X"D3",X"2F",X"B0",X"56",X"DB",X"0D",X"00",X"05",
		X"08",X"A4",X"C0",X"DF",X"FD",X"FF",X"8F",X"3F",X"C0",X"05",X"A0",X"E7",X"5F",X"4A",X"08",X"C1",
		X"14",X"FE",X"05",X"FE",X"DF",X"EF",X"3D",X"E2",X"07",X"00",X"00",X"A0",X"9B",X"5F",X"C7",X"5F",
		X"49",X"54",X"49",X"E1",X"FF",X"77",X"B7",X"FB",X"00",X"E0",X"05",X"80",X"DC",X"03",X"E8",X"57",
		X"26",X"7C",X"87",X"FF",X"FC",X"FE",X"02",X"00",X"FA",X"07",X"60",X"5F",X"04",X"D0",X"7F",X"E0",
		X"F6",X"0F",X"F8",X"81",X"25",X"11",X"F0",X"2A",X"68",X"FF",X"FF",X"A7",X"42",X"04",X"1E",X"8F",
		X"7F",X"4A",X"28",X"E0",X"9F",X"0B",X"1C",X"7F",X"80",X"4F",X"D1",X"07",X"7D",X"E8",X"F6",X"17",
		X"2C",X"00",X"05",X"F0",X"1F",X"FF",X"99",X"FC",X"C3",X"02",X"7E",X"A5",X"EB",X"07",X"8E",X"61",
		X"14",X"80",X"20",X"DD",X"DF",X"FE",X"05",X"21",X"C0",X"87",X"BD",X"F7",X"0F",X"3F",X"04",X"50",
		X"15",X"4B",X"9C",X"7D",X"FD",X"7D",X"AF",X"BA",X"3E",X"58",X"00",X"50",X"1F",X"10",X"44",X"A9",
		X"D4",X"86",X"FF",X"F6",X"5F",X"FF",X"FB",X"40",X"08",X"20",X"F8",X"C1",X"03",X"EF",X"03",X"40",
		X"5E",X"AA",X"12",X"F6",X"7D",X"C5",X"FF",X"47",X"F4",X"07",X"40",X"DE",X"0B",X"80",X"0F",X"FC",
		X"0A",X"89",X"24",X"79",X"D3",X"B5",X"FF",X"17",X"D0",X"FD",X"1F",X"74",X"2F",X"00",X"40",X"57",
		X"EA",X"1F",X"C0",X"3E",X"F0",X"57",X"01",X"EE",X"DF",X"BB",X"9B",X"BC",X"D8",X"02",X"38",X"38",
		X"E0",X"05",X"EF",X"2B",X"25",X"95",X"AA",X"95",X"07",X"F5",X"F5",X"6F",X"D5",X"0F",X"10",X"00",
		X"00",X"C0",X"FB",X"6F",X"77",X"57",X"7D",X"00",X"5F",X"05",X"2E",X"E5",X"E0",X"FF",X"95",X"5A",
		X"55",X"F0",X"DA",X"FF",X"0F",X"1C",X"2E",X"00",X"80",X"6D",X"55",X"D5",X"27",X"00",X"F0",X"13",
		X"11",X"A5",X"60",X"FE",X"FF",X"57",X"EC",X"AD",X"BF",X"80",X"3F",X"70",X"10",X"78",X"78",X"D8",
		X"61",X"F4",X"B0",X"0B",X"20",X"FD",X"DF",X"25",X"F0",X"0D",X"FC",X"8E",X"E3",X"92",X"E0",X"7B",
		X"C6",X"86",X"9F",X"DF",X"41",X"00",X"94",X"D7",X"D7",X"03",X"00",X"55",X"7F",X"0C",X"F2",X"55",
		X"60",X"E7",X"3E",X"09",X"ED",X"FD",X"5E",X"D5",X"1E",X"D0",X"00",X"44",X"12",X"49",X"65",X"0B",
		X"FC",X"FD",X"FF",X"03",X"3F",X"F8",X"80",X"1F",X"38",X"10",X"B0",X"84",X"0B",X"FA",X"FF",X"23",
		X"FD",X"02",X"F8",X"1F",X"91",X"4A",X"8F",X"E0",X"E9",X"81",X"1E",X"FF",X"7D",X"80",X"2F",X"04",
		X"78",X"0B",X"F8",X"F1",X"B0",X"7E",X"14",X"54",X"ED",X"AB",X"7D",X"00",X"02",X"FE",X"98",X"14",
		X"1C",X"FE",X"6B",X"C8",X"BF",X"8B",X"85",X"45",X"C1",X"7F",X"F0",X"A3",X"0F",X"EA",X"32",X"0F",
		X"20",X"01",X"E0",X"F0",X"1F",X"ED",X"3F",X"0B",X"C0",X"FB",X"07",X"BC",X"DF",X"AD",X"9A",X"1E",
		X"00",X"10",X"48",X"51",X"F8",X"FF",X"07",X"FC",X"A9",X"B0",X"67",X"B7",X"81",X"F4",X"03",X"00",
		X"96",X"00",X"7E",X"F7",X"FF",X"C1",X"07",X"E0",X"7F",X"3A",X"45",X"80",X"E4",X"FF",X"A8",X"2F",
		X"7E",X"C0",X"20",X"02",X"67",X"F8",X"FD",X"5F",X"80",X"5E",X"24",X"F0",X"BB",X"64",X"A5",X"0A",
		X"BC",X"7F",X"38",X"08",X"CA",X"EF",X"0A",X"40",X"FB",X"F6",X"5A",X"3F",X"00",X"F0",X"60",X"D7",
		X"BE",X"29",X"80",X"6B",X"F4",X"3F",X"F0",X"B9",X"FF",X"00",X"25",X"20",X"4C",X"04",X"FD",X"C7",
		X"BD",X"B5",X"55",X"0A",X"1A",X"16",X"00",X"12",X"22",X"02",X"FF",X"FF",X"FF",X"C1",X"A3",X"6D",
		X"F5",X"1F",X"40",X"71",X"A8",X"7B",X"01",X"F8",X"A4",X"92",X"14",X"FC",X"FF",X"DA",X"04",X"6A",
		X"59",X"60",X"FE",X"C3",X"2C",X"00",X"AE",X"F5",X"07",X"D8",X"0F",X"E8",X"07",X"03",X"DC",X"0F",
		X"3A",X"7F",X"07",X"40",X"FF",X"3E",X"7C",X"49",X"C4",X"F2",X"55",X"41",X"FF",X"6B",X"7F",X"00",
		X"1C",X"04",X"81",X"FA",X"01",X"8F",X"5D",X"C0",X"FF",X"17",X"F0",X"1F",X"01",X"97",X"0E",X"9F",
		X"AF",X"43",X"68",X"EF",X"C7",X"07",X"4A",X"50",X"70",X"0F",X"BA",X"FF",X"D1",X"FB",X"23",X"24",
		X"70",X"C0",X"94",X"20",X"42",X"05",X"F8",X"FF",X"C3",X"E9",X"1F",X"00",X"3E",X"F8",X"4B",X"80",
		X"5B",X"D1",X"B9",X"B7",X"7F",X"80",X"81",X"1F",X"0D",X"F0",X"1F",X"3C",X"FD",X"61",X"E1",X"07",
		X"CE",X"F5",X"0F",X"01",X"5C",X"FE",X"09",X"F8",X"70",X"28",X"24",X"E1",X"F7",X"C1",X"F3",X"7C",
		X"01",X"7E",X"0D",X"DC",X"D4",X"7F",X"01",X"3C",X"C2",X"63",X"0B",X"95",X"52",X"D8",X"6F",X"FF",
		X"07",X"41",X"70",X"62",X"15",X"D6",X"FF",X"51",X"C0",X"FD",X"CF",X"21",X"3D",X"24",X"80",X"87",
		X"90",X"20",X"3B",X"58",X"5F",X"FF",X"5F",X"02",X"F8",X"FF",X"02",X"BE",X"40",X"47",X"AB",X"DA",
		X"6A",X"59",X"0B",X"0C",X"80",X"7F",X"05",X"FA",X"5F",X"B0",X"BD",X"BF",X"F1",X"31",X"C1",X"00",
		X"9F",X"00",X"A1",X"22",X"AC",X"55",X"F5",X"F7",X"8F",X"04",X"9F",X"E9",X"FE",X"A0",X"FD",X"00",
		X"B0",X"BF",X"00",X"03",X"1F",X"F8",X"FF",X"02",X"FA",X"1F",X"0E",X"BE",X"C5",X"4B",X"C1",X"47",
		X"09",X"FC",X"44",X"FD",X"03",X"5A",X"7D",X"2B",X"C0",X"82",X"50",X"81",X"82",X"EF",X"7F",X"F5",
		X"A5",X"0A",X"0F",X"16",X"25",X"14",X"F8",X"97",X"E8",X"FF",X"CF",X"08",X"96",X"C0",X"0F",X"7B",
		X"ED",X"D1",X"D0",X"7A",X"2E",X"0C",X"78",X"08",X"82",X"04",X"FF",X"DF",X"F2",X"8B",X"E0",X"E1",
		X"5F",X"29",X"5C",X"A4",X"1E",X"5F",X"2D",X"18",X"16",X"C0",X"D3",X"4F",X"E8",X"3F",X"58",X"40",
		X"8A",X"7B",X"D0",X"F7",X"B4",X"8E",X"9B",X"74",X"E0",X"BF",X"4F",X"D5",X"7A",X"C0",X"50",X"D0",
		X"80",X"08",X"29",X"B0",X"BF",X"FF",X"E7",X"45",X"78",X"88",X"F6",X"FE",X"FA",X"00",X"02",X"2E",
		X"6A",X"7F",X"15",X"20",X"55",X"A8",X"F8",X"EB",X"EB",X"76",X"FF",X"05",X"F0",X"84",X"2A",X"09",
		X"78",X"EB",X"02",X"6F",X"F4",X"89",X"AF",X"00",X"BC",X"4F",X"6B",X"37",X"39",X"1F",X"00",X"08",
		X"A8",X"54",X"6B",X"F5",X"68",X"FF",X"DD",X"EF",X"B7",X"2D",X"55",X"01",X"7C",X"80",X"00",X"10",
		X"0F",X"7D",X"7D",X"C1",X"5F",X"4F",X"B5",X"57",X"9F",X"A5",X"1D",X"40",X"E9",X"0B",X"10",X"4C",
		X"44",X"B1",X"AE",X"6B",X"EB",X"F5",X"FF",X"1F",X"14",X"DF",X"00",X"9A",X"84",X"16",X"3E",X"80",
		X"3E",X"21",X"10",X"FF",X"5F",X"13",X"97",X"C2",X"F9",X"3F",X"E8",X"1F",X"EA",X"C3",X"07",X"68",
		X"4F",X"00",X"E0",X"D3",X"0F",X"E0",X"F3",X"05",X"7D",X"31",X"7C",X"50",X"BF",X"54",X"18",X"7C",
		X"C4",X"5F",X"C0",X"2B",X"C1",X"F4",X"4E",X"5F",X"FD",X"30",X"F0",X"F6",X"5F",X"03",X"50",X"49",
		X"00",X"BA",X"BF",X"FD",X"43",X"82",X"4A",X"B0",X"70",X"3B",X"FC",X"FC",X"2D",X"F8",X"80",X"F6",
		X"8F",X"06",X"D0",X"0F",X"1A",X"F1",X"2E",X"F6",X"A7",X"0A",X"F0",X"12",X"1A",X"E8",X"AE",X"7F",
		X"1E",X"65",X"E8",X"40",X"F9",X"03",X"8D",X"EA",X"71",X"81",X"6B",X"0E",X"78",X"F8",X"72",X"F4",
		X"2B",X"A8",X"6B",X"81",X"BF",X"02",X"FC",X"0F",X"68",X"BF",X"A9",X"7E",X"01",X"70",X"05",X"3C",
		X"05",X"DE",X"57",X"E1",X"59",X"7F",X"F0",X"2F",X"7C",X"51",X"A8",X"07",X"BD",X"84",X"3F",X"F0",
		X"42",X"C5",X"8B",X"0F",X"86",X"BF",X"C2",X"08",X"F8",X"81",X"2F",X"65",X"17",X"8E",X"FF",X"1F",
		X"D6",X"05",X"D2",X"31",X"D0",X"71",X"13",X"E0",X"0F",X"7A",X"61",X"BF",X"15",X"E1",X"97",X"40",
		X"F0",X"FD",X"94",X"52",X"5A",X"FD",X"3A",X"3E",X"00",X"AD",X"3F",X"C0",X"07",X"6C",X"5F",X"02",
		X"7B",X"2D",X"D4",X"0F",X"F8",X"07",X"5E",X"45",X"6C",X"7C",X"60",X"51",X"FB",X"D2",X"CB",X"2B",
		X"00",X"FD",X"1B",X"F0",X"1B",X"E0",X"E3",X"3C",X"F0",X"0B",X"B8",X"5C",X"E0",X"E0",X"0F",X"EC",
		X"7F",X"12",X"F0",X"51",X"89",X"EE",X"DA",X"FE",X"28",X"81",X"10",X"C0",X"FD",X"C7",X"5F",X"E0",
		X"2B",X"14",X"68",X"1F",X"3F",X"F0",X"E3",X"80",X"D9",X"6A",X"EB",X"02",X"C3",X"0B",X"00",X"FD",
		X"9F",X"5C",X"D0",X"6F",X"E8",X"2F",X"0E",X"AA",X"08",X"BA",X"E8",X"6B",X"BD",X"76",X"E1",X"43",
		X"18",X"B8",X"70",X"95",X"48",X"60",X"FF",X"F1",X"17",X"7D",X"0B",X"D2",X"A1",X"FD",X"57",X"45",
		X"00",X"50",X"5F",X"82",X"2E",X"BF",X"C7",X"0F",X"28",X"FD",X"8E",X"82",X"75",X"2D",X"A0",X"D5",
		X"FF",X"43",X"13",X"54",X"4A",X"49",X"85",X"FE",X"EE",X"F7",X"17",X"C1",X"0F",X"00",X"F4",X"03",
		X"5C",X"40",X"3F",X"8D",X"7E",X"F8",X"DB",X"04",X"AD",X"12",X"F0",X"6F",X"77",X"FD",X"81",X"0B",
		X"E0",X"02",X"F4",X"8A",X"2A",X"F8",X"83",X"BE",X"FE",X"17",X"29",X"E0",X"2B",X"50",X"FF",X"22",
		X"7E",X"04",X"FA",X"01",X"58",X"5F",X"46",X"EF",X"85",X"05",X"B8",X"68",X"1F",X"4F",X"1F",X"D4",
		X"2F",X"C4",X"57",X"A1",X"58",X"2D",X"E2",X"AF",X"64",X"60",X"AF",X"1F",X"03",X"FC",X"02",X"3E",
		X"60",X"62",X"FF",X"68",X"0B",X"AF",X"05",X"29",X"D2",X"1F",X"EA",X"FE",X"63",X"7F",X"74",X"00",
		X"ED",X"27",X"A1",X"84",X"03",X"7F",X"45",X"E9",X"17",X"28",X"3F",X"C4",X"E5",X"C2",X"0A",X"57",
		X"48",X"75",X"AF",X"4A",X"0B",X"3E",X"68",X"09",X"8E",X"06",X"FE",X"1F",X"57",X"B6",X"02",X"6F",
		X"AF",X"EB",X"83",X"F6",X"81",X"AA",X"EA",X"0E",X"C0",X"17",X"40",X"A2",X"87",X"FA",X"F3",X"B0",
		X"BF",X"08",X"54",X"FB",X"D6",X"27",X"0B",X"7C",X"E4",X"05",X"89",X"3E",X"24",X"FC",X"ED",X"82",
		X"F2",X"75",X"25",X"F0",X"03",X"DA",X"CF",X"E2",X"07",X"45",X"F5",X"41",X"AF",X"80",X"0F",X"BB",
		X"28",X"F4",X"55",X"9A",X"EE",X"E1",X"B7",X"4A",X"95",X"AF",X"20",X"70",X"0B",X"94",X"7E",X"FC",
		X"80",X"76",X"E1",X"03",X"83",X"0F",X"63",X"DA",X"E9",X"2B",X"5D",X"F2",X"34",X"05",X"F6",X"16",
		X"2A",X"80",X"F7",X"7D",X"FF",X"C1",X"01",X"A8",X"1F",X"A0",X"BA",X"3A",X"3D",X"1C",X"2C",X"B0",
		X"F4",X"57",X"16",X"1C",X"F2",X"77",X"45",X"3E",X"F2",X"5A",X"BB",X"14",X"10",X"F8",X"AC",X"EA",
		X"7E",X"A5",X"0A",X"F0",X"95",X"FE",X"22",X"B4",X"1F",X"41",X"22",X"12",X"F8",X"D6",X"5F",X"54",
		X"BD",X"A0",X"FF",X"D0",X"1E",X"16",X"E8",X"12",X"D0",X"03",X"7C",X"D3",X"55",X"35",X"E9",X"43",
		X"E7",X"82",X"A0",X"F4",X"6B",X"4B",X"FF",X"D1",X"02",X"1E",X"54",X"6F",X"81",X"3F",X"42",X"2E",
		X"AF",X"FA",X"25",X"01",X"15",X"3C",X"1D",X"FD",X"93",X"C0",X"EB",X"C3",X"96",X"3A",X"A6",X"AB",
		X"B0",X"80",X"8F",X"57",X"0F",X"D5",X"56",X"55",X"E9",X"FC",X"02",X"79",X"51",X"E8",X"03",X"B6",
		X"7F",X"05",X"A4",X"A9",X"7D",X"81",X"A0",X"51",X"5F",X"92",X"CA",X"E8",X"07",X"FD",X"D7",X"0A",
		X"C1",X"D5",X"BB",X"14",X"81",X"2B",X"E4",X"B2",X"B7",X"D6",X"57",X"10",X"D4",X"AE",X"92",X"80",
		X"3F",X"EC",X"1F",X"1F",X"FC",X"2C",X"57",X"15",X"F4",X"25",X"08",X"5E",X"B1",X"B8",X"2A",X"E0",
		X"D7",X"82",X"5A",X"F7",X"91",X"E5",X"10",X"E0",X"65",X"5F",X"42",X"A9",X"F0",X"FD",X"F2",X"D2",
		X"35",X"05",X"B3",X"D8",X"03",X"16",X"1D",X"F1",X"87",X"5E",X"3C",X"D4",X"0B",X"F4",X"E5",X"B5",
		X"40",X"3F",X"81",X"47",X"43",X"DF",X"AA",X"80",X"F5",X"AA",X"44",X"F2",X"AF",X"74",X"55",X"B8",
		X"0B",X"A4",X"FD",X"05",X"A9",X"97",X"C5",X"A5",X"80",X"E0",X"57",X"AD",X"14",X"FE",X"AA",X"85",
		X"FB",X"2F",X"81",X"EA",X"F8",X"2E",X"B0",X"D4",X"42",X"40",X"7F",X"11",X"56",X"7B",X"94",X"6B",
		X"A1",X"EA",X"45",X"D5",X"D2",X"03",X"DF",X"49",X"51",X"5A",X"09",X"BF",X"FB",X"05",X"DC",X"E2",
		X"15",X"1A",X"55",X"07",X"FF",X"85",X"90",X"AA",X"3A",X"E1",X"7D",X"E0",X"85",X"FE",X"81",X"6B",
		X"A0",X"5F",X"50",X"D5",X"8B",X"A2",X"FD",X"15",X"D0",X"5F",X"82",X"A8",X"5F",X"E8",X"2D",X"78",
		X"9C",X"12",X"E5",X"60",X"2F",X"7A",X"0B",X"B0",X"D5",X"5E",X"95",X"08",X"5A",X"F8",X"86",X"FE",
		X"78",X"D2",X"17",X"70",X"1A",X"95",X"50",X"5D",X"EA",X"FD",X"69",X"05",X"EA",X"81",X"BD",X"82",
		X"17",X"AF",X"F0",X"A8",X"BB",X"B7",X"14",X"98",X"16",X"F0",X"F0",X"AB",X"40",X"7F",X"1B",X"AD",
		X"07",X"D5",X"02",X"C6",X"5D",X"28",X"87",X"7E",X"02",X"57",X"45",X"75",X"6D",X"F8",X"4B",X"6F",
		X"4B",X"3B",X"B4",X"05",X"D1",X"06",X"15",X"01",X"FD",X"46",X"17",X"2F",X"EC",X"7D",X"F4",X"4B",
		X"BB",X"08",X"2A",X"8D",X"02",X"FA",X"5D",X"C2",X"55",X"B2",X"84",X"DE",X"BB",X"AA",X"10",X"9A",
		X"D4",X"17",X"F4",X"72",X"0F",X"07",X"69",X"D1",X"2F",X"94",X"7A",X"58",X"7D",X"05",X"07",X"D8",
		X"BE",X"50",X"5F",X"49",X"E2",X"45",X"55",X"BF",X"F4",X"93",X"40",X"55",X"5D",X"D0",X"B6",X"5E",
		X"14",X"6A",X"07",X"2E",X"54",X"DB",X"E0",X"0B",X"7D",X"45",X"E5",X"9D",X"9E",X"54",X"BD",X"D7",
		X"D4",X"DA",X"01",X"B0",X"5F",X"16",X"A2",X"3E",X"C9",X"82",X"0F",X"5C",X"C5",X"57",X"94",X"AF",
		X"42",X"7D",X"09",X"09",X"FA",X"D5",X"5F",X"08",X"97",X"02",X"F5",X"AF",X"44",X"51",X"A9",X"BA",
		X"17",X"9E",X"58",X"15",X"5C",X"5F",X"89",X"D8",X"57",X"97",X"A4",X"44",X"65",X"4B",X"5F",X"F9",
		X"E0",X"AB",X"45",X"A1",X"78",X"51",X"4B",X"D8",X"B7",X"0F",X"B4",X"8B",X"AA",X"02",X"5D",X"45",
		X"0B",X"55",X"7D",X"BF",X"A0",X"7A",X"69",X"D5",X"15",X"2D",X"0D",X"8A",X"A0",X"3D",X"F5",X"6A",
		X"6F",X"85",X"A2",X"21",X"5D",X"8A",X"2F",X"5D",X"F8",X"F5",X"88",X"2E",X"E8",X"25",X"5E",X"55",
		X"84",X"A4",X"82",X"FB",X"AA",X"F8",X"2A",X"62",X"57",X"5F",X"53",X"41",X"5F",X"45",X"1D",X"1D",
		X"2F",X"A8",X"55",X"04",X"F5",X"17",X"65",X"AD",X"22",X"AB",X"75",X"91",X"5D",X"2B",X"70",X"02",
		X"5A",X"5C",X"47",X"FD",X"55",X"41",X"EB",X"FB",X"40",X"4F",X"54",X"3A",X"F5",X"82",X"94",X"AA",
		X"BE",X"5A",X"A0",X"55",X"75",X"2F",X"70",X"A5",X"22",X"55",X"1F",X"FA",X"FE",X"C5",X"2D",X"54",
		X"B5",X"70",X"95",X"44",X"94",X"EA",X"2F",X"A4",X"56",X"B7",X"D0",X"B3",X"50",X"60",X"AD",X"5B",
		X"48",X"B5",X"AE",X"0A",X"15",X"68",X"FF",X"B8",X"42",X"55",X"55",X"75",X"17",X"54",X"A9",X"6C",
		X"FA",X"0B",X"0A",X"95",X"AA",X"4A",X"85",X"AF",X"DA",X"DB",X"57",X"24",X"C1",X"0A",X"ED",X"EA",
		X"83",X"56",X"D7",X"8A",X"E2",X"A9",X"EA",X"57",X"69",X"41",X"BB",X"17",X"D1",X"17",X"54",X"A5",
		X"BD",X"48",X"75",X"45",X"51",X"5A",X"55",X"C5",X"D7",X"90",X"82",X"56",X"BB",X"EF",X"2A",X"A1",
		X"84",X"9D",X"4A",X"D4",X"4D",X"EF",X"EA",X"A3",X"05",X"55",X"A1",X"D2",X"AA",X"8A",X"9A",X"FA",
		X"82",X"FE",X"1A",X"F4",X"B8",X"52",X"D1",X"A4",X"55",X"AF",X"D0",X"DD",X"28",X"B4",X"A3",X"50",
		X"AD",X"1E",X"D5",X"97",X"B6",X"A0",X"4A",X"BF",X"84",X"B4",X"C4",X"0F",X"55",X"6A",X"85",X"F6",
		X"15",X"FA",X"2A",X"50",X"2B",X"59",X"79",X"74",X"A1",X"6D",X"A5",X"6A",X"BF",X"A0",X"AC",X"82",
		X"2D",X"41",X"FB",X"2B",X"D4",X"A7",X"F6",X"26",X"A4",X"CE",X"85",X"AA",X"17",X"15",X"A1",X"AD",
		X"2E",X"F2",X"55",X"5D",X"45",X"70",X"9D",X"AE",X"56",X"75",X"15",X"21",X"64",X"A7",X"DE",X"52",
		X"08",X"AD",X"8F",X"B4",X"AB",X"EA",X"95",X"28",X"32",X"C4",X"FD",X"57",X"95",X"E0",X"4A",X"A5",
		X"5E",X"55",X"4A",X"A1",X"36",X"81",X"AE",X"A2",X"53",X"B5",X"92",X"FE",X"42",X"AF",X"AA",X"DB",
		X"0A",X"D8",X"2B",X"A0",X"7E",X"49",X"AA",X"D2",X"D7",X"AA",X"C2",X"B3",X"55",X"2B",X"A4",X"2F",
		X"AA",X"22",X"ED",X"57",X"41",X"FA",X"24",X"6A",X"35",X"BD",X"20",X"9A",X"68",X"9D",X"BE",X"84",
		X"D2",X"57",X"7D",X"85",X"AA",X"54",X"5C",X"31",X"8F",X"96",X"5E",X"E8",X"9B",X"50",X"D5",X"A2",
		X"50",X"7D",X"58",X"B4",X"6B",X"1F",X"5D",X"09",X"AD",X"5A",X"60",X"A3",X"CE",X"55",X"4A",X"D5",
		X"4B",X"FB",X"08",X"D5",X"5E",X"71",X"51",X"64",X"A5",X"56",X"92",X"AE",X"2A",X"B6",X"7E",X"05",
		X"56",X"17",X"FA",X"40",X"D8",X"0A",X"0D",X"DA",X"DE",X"BB",X"92",X"2A",X"A5",X"44",X"7D",X"C9",
		X"6B",X"FB",X"A5",X"15",X"D0",X"2F",X"42",X"69",X"55",X"C9",X"F2",X"54",X"D4",X"BB",X"15",X"1E",
		X"52",X"B5",X"2A",X"15",X"DD",X"A4",X"17",X"A6",X"FA",X"B5",X"AA",X"A0",X"5A",X"5F",X"41",X"AF",
		X"12",X"AC",X"15",X"AA",X"55",X"5F",X"21",X"2D",X"4B",X"4A",X"12",X"A9",X"5B",X"6B",X"A5",X"5F",
		X"CB",X"E2",X"2B",X"5B",X"82",X"AA",X"FA",X"10",X"A9",X"2E",X"BD",X"02",X"D5",X"4A",X"A5",X"BA",
		X"55",X"D0",X"AF",X"BE",X"4A",X"45",X"A2",X"BA",X"57",X"B5",X"22",X"97",X"82",X"AA",X"55",X"A1",
		X"6A",X"4A",X"57",X"F1",X"45",X"85",X"AE",X"AE",X"2E",X"B6",X"55",X"91",X"AA",X"76",X"95",X"A0",
		X"AA",X"A4",X"AA",X"FA",X"85",X"2E",X"75",X"15",X"AA",X"5F",X"0D",X"F5",X"15",X"AA",X"AF",X"88",
		X"EC",X"21",X"55",X"D5",X"0D",X"55",X"AB",X"24",X"A1",X"95",X"4A",X"5F",X"61",X"6B",X"DB",X"EB",
		X"2A",X"BB",X"20",X"45",X"8A",X"D4",X"2B",X"F2",X"15",X"FA",X"AA",X"4A",X"55",X"A1",X"97",X"B2",
		X"BA",X"4F",X"A8",X"57",X"A1",X"2A",X"29",X"55",X"55",X"55",X"5C",X"BF",X"96",X"A8",X"AB",X"DA",
		X"57",X"21",X"91",X"A8",X"AA",X"54",X"B5",X"AF",X"56",X"EB",X"42",X"29",X"5D",X"42",X"55",X"B5",
		X"53",X"2A",X"B5",X"AA",X"AA",X"DB",X"25",X"54",X"AD",X"AA",X"52",X"2B",X"B5",X"A2",X"4A",X"91",
		X"52",X"55",X"D5",X"56",X"54",X"69",X"F5",X"A2",X"AA",X"6F",X"A1",X"7A",X"85",X"56",X"15",X"ED",
		X"A0",X"DA",X"95",X"22",X"55",X"A5",X"AB",X"2A",X"55",X"BD",X"52",X"95",X"EA",X"5F",X"85",X"AA",
		X"2A",X"AA",X"0A",X"5D",X"49",X"45",X"D5",X"57",X"A4",X"2B",X"55",X"BD",X"2E",X"AA",X"54",X"A9",
		X"12",X"B5",X"2F",X"AA",X"5E",X"75",X"49",X"55",X"51",X"2F",X"92",X"56",X"2B",X"D5",X"A6",X"A3",
		X"A4",X"56",X"8D",X"5A",X"55",X"55",X"92",X"56",X"AD",X"6C",X"85",X"AA",X"6F",X"AB",X"0A",X"6A",
		X"F5",X"2A",X"85",X"AA",X"AA",X"56",X"AA",X"16",X"D5",X"0A",X"AB",X"88",X"DA",X"DE",X"8A",X"F4",
		X"54",X"F5",X"AA",X"52",X"55",X"A9",X"52",X"55",X"45",X"45",X"95",X"6A",X"AD",X"54",X"B8",X"AA",
		X"AA",X"AA",X"F5",X"5A",X"51",X"2F",X"55",X"AA",X"AA",X"5A",X"55",X"41",X"5A",X"69",X"95",X"D0",
		X"BD",X"A8",X"D6",X"AB",X"56",X"95",X"B4",X"AB",X"95",X"57",X"A4",X"15",X"55",X"55",X"55",X"2B",
		X"55",X"97",X"52",X"D2",X"52",X"15",X"95",X"74",X"55",X"55",X"F5",X"15",X"2A",X"57",X"55",X"AF",
		X"4A",X"54",X"5B",X"A2",X"6A",X"55",X"AA",X"55",X"4B",X"55",X"51",X"AA",X"6A",X"AD",X"AA",X"A0",
		X"4A",X"94",X"5A",X"7F",X"D9",X"55",X"41",X"AB",X"AA",X"56",X"7D",X"45",X"A5",X"AA",X"AA",X"15",
		X"55",X"55",X"55",X"D5",X"4A",X"55",X"AB",X"4A",X"55",X"B5",X"52",X"E5",X"52",X"2B",X"EA",X"57",
		X"A5",X"92",X"4A",X"5D",X"55",X"55",X"A9",X"56",X"69",X"01",X"55",X"ED",X"95",X"54",X"55",X"ED",
		X"A2",X"5E",X"AB",X"15",X"D6",X"AD",X"A4",X"5A",X"55",X"49",X"52",X"AA",X"AA",X"A2",X"AA",X"FA",
		X"54",X"25",X"55",X"55",X"5D",X"55",X"2A",X"BA",X"54",X"2F",X"7A",X"A5",X"52",X"A5",X"56",X"EA",
		X"EA",X"AA",X"52",X"A5",X"5A",X"15",X"55",X"2B",X"6A",X"D1",X"2A",X"5D",X"97",X"94",X"AA",X"55",
		X"A5",X"55",X"F5",X"48",X"AD",X"54",X"B5",X"4A",X"54",X"57",X"A9",X"A4",X"56",X"A9",X"56",X"55",
		X"D5",X"FE",X"52",X"AD",X"BA",X"92",X"48",X"55",X"55",X"45",X"5A",X"55",X"D5",X"9D",X"A2",X"D5",
		X"AA",X"57",X"A5",X"4A",X"25",X"55",X"95",X"52",X"55",X"15",X"55",X"F7",X"55",X"52",X"95",X"EA",
		X"4A",X"55",X"F5",X"AD",X"22",X"55",X"55",X"55",X"D5",X"96",X"A8",X"AA",X"DA",X"2A",X"55",X"A9",
		X"AA",X"6A",X"55",X"55",X"95",X"AA",X"D6",X"AA",X"AE",X"54",X"29",X"52",X"55",X"57",X"A9",X"55",
		X"15",X"29",X"55",X"AF",X"AA",X"92",X"AA",X"AA",X"A8",X"6D",X"AB",X"92",X"54",X"AB",X"2A",X"AA",
		X"56",X"D5",X"AA",X"52",X"55",X"09",X"55",X"55",X"D5",X"AB",X"AA",X"D6",X"45",X"A9",X"ED",X"15",
		X"D5",X"4A",X"A8",X"56",X"25",X"55",X"B5",X"6A",X"55",X"55",X"95",X"AA",X"94",X"AA",X"55",X"A5",
		X"AA",X"6B",X"ED",X"45",X"D5",X"AA",X"44",X"A9",X"4A",X"B5",X"AA",X"AA",X"6F",X"57",X"54",X"A5",
		X"A5",X"AA",X"AA",X"A8",X"6A",X"AD",X"AA",X"68",X"55",X"51",X"D5",X"5A",X"15",X"55",X"D5",X"55",
		X"5F",X"51",X"55",X"95",X"A4",X"BA",X"92",X"AA",X"55",X"A5",X"AA",X"B5",X"56",X"55",X"55",X"44",
		X"55",X"55",X"55",X"AD",X"AA",X"55",X"B5",X"2A",X"AA",X"AA",X"5A",X"6D",X"15",X"AA",X"4A",X"55",
		X"B5",X"AA",X"AA",X"55",X"D5",X"AA",X"A4",X"2E",X"AA",X"6A",X"55",X"55",X"A9",X"8A",X"AA",X"55",
		X"DA",X"AA",X"5A",X"D5",X"92",X"AA",X"AA",X"4A",X"55",X"55",X"D5",X"55",X"A5",X"BA",X"95",X"AA",
		X"AA",X"4A",X"55",X"55",X"AD",X"4A",X"55",X"55",X"54",X"A5",X"AA",X"6A",X"55",X"55",X"55",X"55",
		X"A1",X"AA",X"54",X"55",X"5B",X"AB",X"2A",X"55",X"55",X"55",X"B5",X"2A",X"55",X"A5",X"54",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"B5",X"AA",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"55",X"55",
		X"B5",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"55",X"55",X"55",X"A9",X"AA",X"AA",X"AA",X"AA",X"54",
		X"55",X"55",X"55",X"55",X"55",X"D5",X"AA",X"AA",X"AA",X"AA",X"54",X"45",X"55",X"55",X"55",X"55",
		X"A9",X"AA",X"AA",X"AA",X"AA",X"52",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A9",X"AA",
		X"AA",X"AA",X"6A",X"55",X"55",X"55",X"51",X"45",X"55",X"55",X"75",X"55",X"A9",X"BA",X"AA",X"AA",
		X"AA",X"AA",X"4A",X"55",X"55",X"AD",X"AA",X"4A",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"AB",X"AA",X"5A",X"55",X"55",X"55",X"95",X"AA",X"52",X"55",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"B5",X"AA",X"AA",X"5A",X"55",X"55",X"55",X"55",X"55",X"55",X"A9",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"55",X"AA",X"AA",X"AA",X"6A",X"55",X"55",X"55",
		X"55",X"55",X"55",X"A9",X"AA",X"52",X"55",X"55",X"55",X"55",X"55",X"AD",X"AA",X"56",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A5",X"AA",X"AA",X"AA",X"AA",X"2A",X"55",X"AB",X"AA",
		X"AA",X"AA",X"54",X"55",X"55",X"95",X"54",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"A9",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"5A",X"55",X"55",X"55",X"55",X"95",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"54",X"55",X"55",X"55",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3B",
		X"4F",X"C6",X"00",X"F7",X"78",X"00",X"20",X"FB",X"86",X"01",X"20",X"F5",X"86",X"02",X"20",X"F1",
		X"FF",X"E8",X"FF",X"E8",X"FF",X"E8",X"FF",X"E0",X"FF",X"E8",X"FF",X"E8",X"FF",X"EC",X"FF",X"E8");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
